 library ieee;
 use ieee.std_logic_1164.all;
 use ieee.numeric_std.all;
 
 entity ram_l1_n4 is
	generic(
		g_width 		: natural := 16;
		g_depth 		: natural := 50;
		g_addr_bits : natural := 5);
	
	port(
		i_clk			: in std_logic;
		i_wr			: in std_logic;
		i_addr		: in std_logic_vector(g_addr_bits-1 downto 0);
		i_data		: in std_logic_vector(g_width-1 downto 0);
		o_data		: out std_logic_vector(g_width-1 downto 0));
 end ram_l1_n4;
 
 architecture rtl of ram_l1_n4 is
	type t_mem is array (0 to g_depth-1) of std_logic_vector(g_width-1 downto 0);
	signal r_mem 	: t_mem := ("1110110011111001", "0000000010111000", "1111110011100101",
									 	"0000001010001011", "0000010001000101", "1111111101111100", others => (others=>'0'));

 begin
	p_ram : process(i_clk)
	begin
		if rising_edge(i_clk) then
			if (i_wr='1') then
				r_mem(to_integer(unsigned(i_addr))) <= i_data;
			end if;
			o_data <= r_mem(to_integer(unsigned(i_addr)));
		end if;
	end process p_ram; 
 end rtl;