library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram_l4_n3 is
	generic(
		g_width   : natural := 16;
		g_depth 	: natural := 50;
		g_addr_bits : natural := 5);
	port(
		i_clk			: in std_logic;
		i_wr			: in std_logic;
		i_addr		: in std_logic_vector(g_addr_bits-1 downto 0);
		i_data		: in std_logic_vector(g_width-1 downto 0);
		o_data		: out std_logic_vector(g_width-1 downto 0));
end ram_l4_n3;

architecture rtl of ram_l4_n3 is
	type t_mem is array (0 to g_depth-1) of std_logic_vector(g_width-1 downto 0);
	signal r_mem : t_mem := ("0000010011011100", "0000101010010001", "1111110110011110", "1111101011100011", "0000110011100110", "0000000111000110", "0000010000011111", "0000000001110111", "1111010000011011", "0000001100001111", "0000001000001001", "1111101010010010", "0000010111100001", "1111111000010110", "0000011110101010", "1111010100000000", "0001010001001100", "0000010000110110", "1111101110100011", "0000001110011101" , others => (others => '0'));

begin
	p_ram : process(i_clk)
	begin
		if rising_edge(i_clk) then
			if (i_wr='1') then
				r_mem(to_integer(unsigned(i_addr))) <= i_data;
			end if;
			o_data <= r_mem(to_integer(unsigned(i_addr)));
		end if;	end process p_ram;end rtl;