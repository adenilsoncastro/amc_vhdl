library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram_l4_n0 is
	generic(
		g_width   : natural := 16;
		g_depth 	: natural := 50;
		g_addr_bits : natural := 5);
	port(
		i_clk			: in std_logic;
		i_wr			: in std_logic;
		i_addr		: in std_logic_vector(g_addr_bits-1 downto 0);
		i_data		: in std_logic_vector(g_width-1 downto 0);
		o_data		: out std_logic_vector(g_width-1 downto 0));
end ram_l4_n0;

architecture rtl of ram_l4_n0 is
	type t_mem is array (0 to g_depth-1) of std_logic_vector(g_width-1 downto 0);
	signal r_mem : t_mem := ("0000011111001111", "0000001100000100", "0001000110011111", "1111111100101010", "0000011110011100", "1111111111111001", "1111111101111010", "0000010011000101", "1111011010010000", "0000000000010001", "1111000110000110", "0000011101111010", "1111011001000011", "1111011100010011", "0000010010011011", "0000000010011111", "1111110100101000", "0001000101101010", "1111111111011110", "0000111110111011" , others => (others => '0'));

begin
	p_ram : process(i_clk)
	begin
		if rising_edge(i_clk) then
			if (i_wr='1') then
				r_mem(to_integer(unsigned(i_addr))) <= i_data;
			end if;
			o_data <= r_mem(to_integer(unsigned(i_addr)));
		end if;	end process p_ram;end rtl;