library ieee;
use ieee.std_logic_1164.all;

package data_types is
	type complex is record
		re		: std_logic_vector(15 downto 0);
		img	: std_logic_vector(15 downto 0);
	end record;
	
	type mod_data is array (0 to 5) of complex;
end data_types;
