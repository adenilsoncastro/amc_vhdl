 library ieee;
 use ieee.std_logic_1164.all;
 --use ieee.numeric_std.all;
 
 library ieee_proposed;
 use ieee_proposed.fixed_pkg.all;
 
 library rna_library;
 use rna_library.data_types_pkg.all;
 
 entity features is 
	generic(
		g_bits			: natural := c_bits;
		g_fxp_high		: natural := c_fxp_high;
		g_fxp_low		: integer := c_fxp_low;
		g_frame_size	: natural := c_frame_size);	
	port(
		i_clk		: in std_logic;
		i_rst		: in std_logic;
		i_enable	: in std_logic;
		i_input 	: in std_logic_vector(g_bits-1 downto 0);
		o_ft_0	: out std_logic_vector(g_bits-1 downto 0);
		o_ft_1	: out std_logic_vector(g_bits-1 downto 0);
		o_ft_2	: out std_logic_vector(g_bits-1 downto 0);
		o_ft_3	: out std_logic_vector(g_bits-1 downto 0);
		o_ft_4	: out std_logic_vector(g_bits-1 downto 0);
		o_ft_5	: out std_logic_vector(g_bits-1 downto 0);
		o_done	: out std_logic);
 end features;
 
 architecture bhv of features is
 
	-- ABS/Mean/
	signal r_ft_state : std_logic_vector(7 downto 0) := (others => '0');
 
	-- Memory arrays
	type t_mem_real is array (0 to g_frame_size-1) of std_logic_vector(g_bits-1 downto 0);
	type t_mem_img is array (0 to g_frame_size-1) of std_logic_vector(g_bits-1 downto 0);
	type t_mem_abs is array (0 to g_frame_size-1) of std_logic_vector(g_bits-1 downto 0);
	type t_mem_cn_abs is array (0 to g_frame_size-1) of std_logic_vector(g_bits-1 downto 0);
	
	signal r_mem_real 	: t_mem_real 	:= ("0000000110010011","1111101101101001","1111110101111100","0000000110110001","1111100011100110","1111110011000101","1111100001101001","1111101100001100","0000001110101001","1111011010011000","1111101101100110","1111111000010001","1111011000011101","1111111101011001","1111001100011000","1111111100100101","0000000010011111","1111011111100100","1111110010011000","0000001011110000","1111111011001111","1111011011001111","0000000101101101","0000001100000010","0000000111110000","0000001111100001","0000001110011101","0000011111111110","1111101011101011","1111011001110011","0000001111101001","1111110100111011","1111011111110111","0000010000001100","1111101100000010","0000001001011000","1111111101110100","0000010101000110","0000000000001101","0000000101110000","1111101100010000","1111101111000000","0000100000110111","1111111001001000","0000000110011001","1111100001100010","0000010010100011","0000000011111001","0000001111111001","0000000000011100","1111101100111010","0000100110011100","0000000011110101","1111010001001101","0000000000010001","1111101101101001","1111111001101111","0000011001011001","1111110000110110","0000011111101011","0000000101001111","1111101000001000","0000101011101100","0000010001111010","0000010100110001","1111101000110100","0000011011101110","0000010110010101","1111110110000010","0000011010010101","0000010011011011","0000010001101011","0000010011111010","1111110100110010","1111100110010110","1111110000111001","1111011111101011","1111110101010100","0000001110011011","1111111100111000","0000000000111000","0000001010010110","1111100111101011","1111110001101101","1111111110111000","0000010101001000","1111111100101111","1111001100000110","0000001001001101","1111100011110111","0000010001011110","1111110011110000","0000011010011001","0000001001100001","1111111101110010","1111100101110110","1111101001000000","1111001101110011","1111000111000001","1111010101111110","1111100100111101","1111111110010111","1111111110001011","1111100111110101","1111100011111011","0000010100000111","1111111101100111","1111110001111011","1111110001010011","0000000100100110","1111010111001100","1111111111011111","0000000110010001","0000010111110111","1111101011111001","1111111000010000","0000001000100110","0000011010101101","1111011001011100","1111010010110001","1111101111010101","1111111001110000","0000000110011011","0000000011011110","1111110100110000","0000010011101101","0000000111110111","1111111101111001","0000001000100100","0000100001011010","0000010000000010","1111111011011101","1111011011110001","1111111010100011","0000000001111111","1111110010101101","0000000100000110","1111100000010010","1111101111010111","0000000001100111","1111010010010111","1111111111110111","1111111000110111","0000010111110101","1111101100110011","1111010110100110","0000001110000001","0000011000000011","0000010011010111","0000101000001100","1111101000111111","1111110000100101","0000010001010011","0000100000010000","0000110111001100","0000000100010100","0000000101010000","0000001100111001","1111110101000000","1111111000101000","1111111010101101","1111111100001010","0000100010011011","0000010100011000","1111110111100101","0000001100010110","1111110010101011","1111111011010110","1111101001110010","0000000111110000","1111101000011001","0000111101001110","0000010011101101","1111100000001011","1111110001101100","1111101110111001","1111010001100010","0000001100100110","1111101111011011","0000010000000001","0000000001010110","0000001011001111","0000000001011110","0000101111001110","1111111000111111","1111111101101100","0000010000000000","1111110001111011","1111110111100010","1111111101001101","1110111100110111","1111111100001010","1111110101101110","0000011001101001","1111110011110100","0000100011110101","0000000110011101","1111110101111111","0000011010000111","0000001001001010","1111111111000101","0000000100101001","0000010000001111","0000100010010000","1111111100001010","0000001110010000","0000000001011100","0000001001100100","1111111101110100","1111111111000000","1111100101010101","1111111101110010","1111111110001000","1111111111011011","0000001111100000","0000001110100101","1111111111000000","1111110011010011","0000001000001110","1111111100000100","1111111010110010","0000000000000000","1111111100010010","1111111101101110","0000001110010000","0000000011111101","0000100100010001","0000010110110101","1111111001111010","0000000111101101","0000000001010011","0000001110000001","0000110010011111","0000101001011010","0000001101111110","1111111101001010","1111110010101110","0000010110010100","1111111111000010","0000000111100101","1111111100001011","1111111110111011","1111111001111011","1111111101010010","1111111010011111","1111110101100000","1111101100111111","1111010010110010","1111101111110001","1111100110111000","0000000110011101","1111101011001010","0000011010111000","0000000110000001","0000001001110111","1111111101100100","1111100011001010","1111110101111110","1111101111000110","1111011101011001","0000000001010011","1111110001001101","0000010101001110","0000010011000000","1111101111000001","1111100011000100","1111101000101110","1111111110001101","0000000011010011","1111101110010101","1111101111010001","0000001110010000","0000000010111000","0000001111110000","1111111001100110","1111011101101110","0000001001001100","0000000110011001","1111110111111110","0000010000010001","0000000111100011","0000001111101010","1111010010010000","0000001110011010","1111111101111001","0000000111000111","0000011101010011","1111101100110101","1111111011111110","0000010001111001","0000011010001010","0000000111101111","0000011010111011","0000100000010010","0000011001111000","1111111100011110","0000010010100011","0000010110101010","0000001010000100","0000011011000100","1111011110111111","0000100010011110","0000001001100111","1111101111100000","1111101111011111","0000000011100011","1111101001101110","0000001010101100","1111110010001011","1111111101000100","0000010101001101","1111011110001000","1111100101011010","0000010111101010","0000000000010100","0000111101001000","0000001000100000","0000000111000101","1111101111000001","1111110111100000","1111100110001101","1111101101100000","0000011111110001","1111101001101111","1111110100101100","0000011111100111","0000001000000010","0000000110011111","1111011010101001","1111110101001010","1111111101111111","0000011011010101","1111101110110001","1111110100010100","1111101111101100","0000100000101000","0000000100101011","1111011001111001","0000001001110000","1111110001010100","0000011001001000","1111111100000010","1111110011111001","0000001010001011","0000010011100110","1111111100011000","0000011001011010","0000000010000000","0000000000110111","0000100100110101","0000001010010110","1111011001010011","0000000001010001","1111110111001000","0000000110101101","1111100110100101","1111100110011101","1111011111101100","1111110110011011","1111010101101010","1111111110000000","0000001100000100","0000000110011001","0000010000001001","1111100111010010","0000001001001100","1111110001000010","0000010001100111","1111111010110001","1111011011101110","1111011101000110","1111010111110100","1111100001110001","0000000000100110","1111101111110111","1111001011111110","0000101011101011","0000000000110011","0000011101110001","1111111101000101","1111111101101001","1111111100111100","1111111011011010","0000100111001000","1111101111110001","0000110111011000","1111010011010000","1111111110001100","1111011001001000","0000000011011000","1111010110001010","1111111100100101","1111100010110110","0000100110001010","0000001110011010","0000011100100010","1111101110000100","1111011101111100","1111011000101001","0000000001011010","0000010100111011","0000101011100111","0000001110101111","0000001010011100","0001000110111101","1111111101100100","1111110011010101","1111110010010011","1111011111011001","0000100110110101","1111100001100110","1111101111111000","0000010110100101","1111110011010000","0001000010000110","1111111011010011","1111100111111001","0000000111100111","1111101011011110","1111111011000000","1111111111110010","0000101101000011","1111101100000010","0000010100010001","0000100101110100","1111110101101011","0000000111110100","1111110010101100","0000101000111010","0000000100001100","0000000110110101","1111110110001000","0000000001011011","1111101100000110","1111000001111000","1111111001100101","1111100100100100","1111111000111001","0000010100011100","1111110110100000","1111011100011011","1111111000100111","0000101010111000","0000011110010101","0000010011111000","0000100010000110","1111111001001001","1111101011101110","1111110110010111","1111111111101000","1111100111000000","0000001011111101","1111111110010011","0000010101011001","1111110100111010","0000001111011110","1111101011001110","0000001001100111","1111111010001111","1111101011011011","1111111000011011","0000000011110000","1111111011110101","1111111011100010","1111100010000011","0000000001000100","1111111100010010","0000010001000100","0000011100011001","0000000000011000","1111010010011100","1111101000110001","1111101110000101","1111110101101000","1111110100001100","0000011101111010","1111010001100100","0000010110011001","0000000101001000","0000000110010111","0000000011011001","1111111101111010","1111111000011111","1110111000001100","1111101101011001","1111111010100110","0000001011110101","1111111001001001","1111110111100111","1111100111001011","1111101000110100","0000000110001101","1111011011101001","0000001010110101","1111100101101111","1111101011100111","1111111001100110","0000000110110010","1111111001000010","1111110001001001","1111111110001101","0000000100000101","0000010111010100","0000010101101101","1111110001011000","1111010110010001","0000000111100010","0000010110111010","1111000000100110","0000001101000001","0000001100110111","1111110110110110","0000001000001011","0000000101011111","1111100111010000","0000010001011101","0000010001100011","0000000010101111","0000001010100100","1111111110011100","1111101101010100","0000000000100100","0000000110100010","1111110011000000","1111111110011101","1111101010011000","0000000100001000","1111101000110001","0000000110011000","1111110101010001","0000001101011010","1111111010010110","1111100011101001","0000010010101000","1111101010011110","0000001011101100","0000010000010110","1111111011111001","1111110011111101","1111111000111111","1111101111111100","1111111100011110","1111110010101101","1111011010010010","0000010011010100","0000011101110001","1111110100010101","1111101111100000","1111101111110000","0000100110011001","0000010100001101","0000000111101101","1111111001101111","0000011100001010","0000000001011110","0000010100001010","0000001010100010","0000000101011111","1111110000101011","0000110000100111","1111110001101110","1111100011010011","0000000001001111","0000000000000011","1111110011000111","0000010010100101","1111111110001010","0000001110111001","0000100001100001","1111100111100111","0000001111011011","0000100101000000","0000001101010110","0000010001011101","0000000001100000","0000010011100001","0000010011101110","1111111101111110","0000010101010110","1111011100111000","0000100010011100","1111110001010001","0000000001011111","1111111100001011","1111111000101100","0000110000110110","1111111011100101","0000001001010101","0000000111110011","1111111000111011","1111110000000111","1111011110100010","0000000111110011","1111110011101011","1111110011101000","1111010110101000","0000010010111100","1111010111100010","0000100101111001","1111001011110001","1111111110011001","1111000110010111","0000000011011110","1111101000011100","0000000010100011","0000010001000110","1111110100101100","0000001010001111","1111110011110000","0000100000101011","0000011010101000","1111110011101100","0000110010110000","1111000110111000","0000001110101110","1111111110011001","1111110000111110","0000000011111001","0000001100010101","0000111101010100","1111110000011001","0000010000101011","0000011001001100","0000000110100100","0000001011110110","0000100001010110","0000000001011101","0000010011111111","0000011100111110","0000001111101100","0000000001100010","0000001010111000","1111011011101111","0000010100000000","0000100110010110","1111110011010001","1111111001010000","1111110110011010","1111110000101110","0000010110011011","0000001000100101","1111111101011001","1111111001011111","1111110101111100","0000010011011100","0000000001001101","0000000010100011","0000000011110000","0000011101110011","0000000000101010","1111111110000101","0000001111011110","1111111000101101","0000000011110101","1111111100010010","0000010001010011","0000100000011100","0000000001110001","0000010101110111","0000000000111100","0000010011110000","1111110001111001","1111111010111110","0000001011111010","0000000100111011","0000011110110110","1111111000001010","1111110110101100","0000001100101100","1111010100000101","1111111110000111","0000101010000000","1111111010011001","1111110000110000","0000011011101011","1111100000100000","0000010000001010","0000001000011001","0000110010000011","0000010000000100","0000010100000110","1111100000110001","0000100111100100","1111111000000001","1111110111000101","0000101101001110","0000010011111110","1111110111100001","1111100001001110","0000001111000001","1111110101011101","1111010010011010","0000011010111111","0000001011010000","1111110110100101","0000010100010000","1111110011111110","0000000001010000","1111111000010000","0000000000100101","1111100001000001","0000111010011000","1111111011110001","1111101001100110","1111111000110011","1111011101000011","0000001101001001","0000000100001100","0000000010010111","0000100000000000","0000000011101110","0000001010010100","1111110110101111","0000000100000010","1111101011000100","1111101100110101","1111001101011010","1111101011100101","1111011100110000","1111110001011010","0000001000111000","1111110100111111","0000011011001001","0000001001111010","1111111100101001","0000010110000011","0000001101100100","1111111000001010","0000011111011100","0000000100110001","1111111001011011","1111111110101000","0000000101011111","1111110010110001","0000010010011110","1111110100000001","1111111101111111","1111111000111111","0000001101000000","0000011111110110","1111011000101111","0000000011011001","0000011101110000","0000000000011000","0000100001101011","1111111010011100","0000010110001101","0000010100110100","0000000011100001","1111110010101010","0000000011110100","0000011101110100","1111111010111100","0000011100100110","1111011110001100","1111110001101101","1111100100101110","0000000101000101","0000000111001001","0000001010101010","1111110100100101","0000000110101110","1111101000100111","1111110111010000","1111111001000111","1111110101000000","1111101101110100","0000001001011011","0000010010001100","0000001111010001","0000001110110000","1111110010001100","1111101000100100","0000001001101110","0000101010001110","1111011011011010","0000000001011101","0000000000011011","0000000010011000","1111100110001000","1111110000000100","1111100110000110","0000010100011110","0000010011000001","1111110101001100","1111111010111010","1111011011001111","1111111001010111","1111110000001100","0000011101010110","0000001001100001","0000000100111100","1111101111111001","1111111010000001","0000111110001001","0000011100000101","1111111011111101","0000000100000001","1111111110110111","1111110110011011","1111110100000110","1111111100010011","0000001011101001","0000001010000010","1111111110011111","0000010000010101","1111011101101001","0000000111111101","1111010110010101","1111110011101011","1111101101011100","0000000011000010","1111001000001101","1111101000110111","1111010110011111","0000000010100000","1111111110100010","1111110101111001","1111110101101001","0000010100101100","1111111001111111","1111111100110010","1111101100011011","1111111101010100","1111110110011001","1111110110000000","1111110000100110","1111110100000001","1111110101101111","0000010100010011","1111101100000111","0000001101011010","1111111111011010","0000011010001101","1111110110011001","1111101111100001","0000011100110100","1111000111110011","1111111000101000","0001000001010111","0000000111100111","1111011001101100","0000000101111100","0000001011000000","0000010010000000","0000011101011011","1111111001100010","0000000111100101","0000000110011000","1111110111111101","1111111000001111","1111100010010100","1111101010011010","1111011111010001","1111111101001100","1111110110101001","1111110101110110","0000011011101011","0000000001000001","1111111111100001","1111110111000011","1111011111011100","1111111101101110","1111010011110011","1111111010010011","0000000101111100","0000011111010001","1111110000101001","0000000110100110","1111111101110001","1111001011011101","1111010010000110","1111110101001001","0000010011100111","1111101100111111","0000001001111111","1111101101110001","1111101000101001","1111100110001010","1111111111100101","1111111000011010","0000010000010111","1111101010000011","1111110100101101","1111101111011011","1111110010001001","0000010101110111","1111111101011011","1111111001101110","0000000111000100","0000011000011010","0000101010010110","0000100000100101","0000011010101000","1111010011110111","1111010101110110","1111111000100000","1111101010000010","0000010000110010","1111111000000011","1111111011110101","0000001100100011","1111111000010110","0000000111000011","1111101110100111","1111101101001111","1111101011010110","1111111100001100","1111100110101110","0000001001110011","1111000011011010","1111101110010111","0000000101001111","1111101110010011","1111110101011100","0000000000011100","0000000010010011","1111101010000111","0000001110011010","0000101100001011","0000011000010110","1111111001101001","0000001010001001","1111111100010011","0000001001010001","0000101111011011","1111111001101110","0000011000100110","1111101110011110","0000001011001100","1111111010101010","0000010010100100","0000010110111010","0000010010100000","0000000110100010","1111110001011000","1111001111100101","1111111011111000","1111100100010100","0000010100110111","0000000110010000","1111110110011100","0000000100101110","1111111011000000","1111001110100011","1111110000111001","1111100011100011","1111101110101011","1111010101011010","0000001000111010","0000000101100010","0000001010110100","0000000001111001","0000101010110101","0000000001011000","1111100111001011","0000010100111111","0000001111101101","0000001101000010","0000001001001101","1111011101100010","1111100110000011","1111101010101001","1111110001010110","0000001000101010","1111011010101101","1111110101111110","1111001001011101","0000001100110011","0000001001101111","1111100011111001","1111111110100100","1111110001101011","0000111010111101","0001000000001010","0000010010110000","0000101101011101","0000000011100010","0000011110101100","1111111111011110","1111101101010101","0000101001000100","0000001110110100","1111101000101010","0000100011010111","0000010100101110","0000001100111010","0000001010001100","1111110111001001","0000001100001011","0000100001001011","1111101000010100","1111100100110001","0000011110001000","0000001101101111","0000000101001110","1111101111000000","1111100101011000","0000001111111110","1111110100000000","1111011100001010","0000000100101001","1111101001000010","0000010000110101","0000010101111110","1111111000010011","1111111110111101","1111111010011100","0000000010100000","0000001001010110","1111100111111100","0000010010000011","1111111110101010","1111011101001111","1111100101100001","0000000010101010","1111011110000111","1111100100011011","1111100011011001","0000011010101011","0000000010101010","0000001100110100","1111101100101000","1111111110101000","0000000000111111","0000000011000010","1111100101110110","0000010101001110","0000011110000110","0000000011100000","1111101011101101","0000011001001001","1111101000001011","1111111100110010","0000011000111000","0000001110101100","0000101110110010","0000001001101111","0000100010000011","0000011010000111","1111110001110001","1111111001100011","0000001010111110","0000000001001111","1111011001110001","0000010001110001","1111110001001100","1111101000111010","0000011101100010","1111100000110010","1111110010110000","1111001110110010","0000100100001011","0000000111001000","1111110110010010","0000010111001110","0000000101101010","0000000001101100","0000010000100001","1111111000000000","1111110010001110","1111111011010100","0000000001000011","0000010011011000","0000001110100111","1111101011100001","0000110010100101","0000010000011001","0000001000101110","0000001000010111","1111011110011110","1111110110110101","1111110100001011","0000000010001011","1111111000100000","0000000101010100","0000001100111111","0000010010010001","0000001011000010","1111010000011111","0000010001100011","0000011110110011","0000100100110000","1111101010001010","1111100111101011","1111110011111000","1111101110010100","0000010001100011","1111111110010110","0000001001011101","1111111000101011","1111100100000001","1111001111000001","1111110101010101","1111100001000001","0000010110111111","0000001111011000","0000010101100110","0000000110010011","1111110100100111","1111110101001111","1111111101100101","1111101101001010","1111011100010110","0000010000100111","0000001100100101","1111101010110101","0000000100011010","1111110000011000","0000010111111110","0000000001011000","0000000000101010","1111101000110010","1111111111000111","0000000111101000","1111110010011100","0000100111001101","0000101011100010","1111110100011111","0000010001101001","0000101100100010","1111101011001111","0000101100101011","1111101011110011","0000011011110001","0000001100000000","1111111011100101","1111111010110101","0000010011101100","0000001110101000","0000100101101001","0000001110000011","0000111011001011","0000010000011001","1111101000100000","0000000100111101","1111110110010011","0000110010111010","1111111010011011","0000110001111010","0000000000101110","1111110001101101","1111100001110010","1111101100011000","1111001011001111","0000000010010110","1111110110010111","0000101011111101","0000110001011001","1111110000111100","1111111110100000","0000000010110110","0000001001110011","0000010001010011","0000001000001001","0000000101101011","0000000010011010","0000101001101011","1111100010111110","0000011111101010","1111110100000001","0000011100001001","1111111011101101","0000011111000101","1111101010100011","1111011101000000","0000001100000010","1111111011001101","1111110010000000","1111100100101100","1111100011000010","0000001100001001","0000100001111101","0000001100010001","0000000011101111","0000110010101011","0000000110111011","0000000000111101","1111111010111001","0000111111001100","1111110111100110","1111111111000111","1111111001000000","0000010100001000","1111110001110000","1111101110110101","0000000100111100","1111101101000001","1111101000110111","0000010100011001","0000001110010111","1111111111011000","1111101101011100","0000000110111000","0000000111100110","1111101101101000","1111100010110111","0000101100101111","1111110101001000","0000001101100010","1111011111011110","0000000110001011","1111111001010010","1111111010110001","1111101000111110","1111110001100001","0000001110010111","0000001100011111","0000011110111100","1111010010100010","0000011010100100","0000000011101100","1111101101100101","1111110101101101","1111101011011101","0000010111111110","0000000111101010","0000010001101001","1111101110111111","0000001000011000","1111111011010010","0000010000101110","1111110111111011","0000000011000000","0000001000000000","1111101111100000","1111111100011110","1111110100110011","0000000011000011","0000010001001101","1111110110111001","1111101110001000","0000011101101001","1111111110011111","1111110000101101","0000000001010010","1111110100101011","1111100100001011","1111110011100000","1111110010110111","1111100101000011","0000010111100001","0000000110100011","0000000101011111","0000010010011000","0000000111001100","0000010001101111","0000101010111000","0000101100011111","1111101011011000","1111101000111010","1111101101110010","0000001010000110","1111011000110111","1111010100111000","1111111001110100","1111001101011110","1111110000110001","1111111100010111","1111111000101000","0000000000111101","0000000011010110","1111111010010100","0000010100010001","0000010010011110","0000001111101010","0000001010011011","1111111111011011","0000010001010000","0000101011111100","0000001110011010","0000101000000010","0000000000100100","0000001111001101","1111110010101000","0000001010100100","0000000110001101","1111000100010110","0000000111100110","0000011101001000","1111100111111010","0000001011000010","0000011000011101","0000010011011000","0000010011111100","1111011111110010","1111110110011001","0000011011010100","0000100010110111","0000001100000001","0000100011111111","0000100101000010","0000110000000110","0000110111001001","1111001110011010","1111101100111011","1111110101100011","0000011010011011","1111110001111001","0000010110000011","0000010101111011","1111111110000110","1111110101001011","1111110001100100","1111110010101011","0000010110101111","0000001100011111","1111100101100100","1111010000011111","0000011110010010","0000001000101000","1111110010010010","0000010111010111","1111110111111111","1111110110101100","0000101001001001","0000100111001000","0000000010101110","0000011100111111","0000101101001011","0000000110101101","0000000000000101","0000010111001101","0000000110110101","0000010010011001","0000101011011100","0000100000010001","1111111011100011","1111000101101110","1111110110011000","0000000100110011","1111110111010001","0000001011100001","0000011100001101","1111101000111101","0000100010001111","0000100100111110","0000101111101111","1111011100011010","1111100101110101","1111001000001100","1111110101010010","1111100111011110","1111111100001000","1111110110101100","0000101011100010","0000000111111100","1111111001110010","0000001010100010","0000011010111100","1111110010000111","0000011000001100","0000100111010101","0000001010011000","0000100110111010","1111110001010011","1111111001110111","1111001111100000","1111110000111110","0000011001111010","1111101011101100","0000011000011010","0000010110101100","0000100000010110","1111100001100001","0000011000001101","0000001100001000","1111110001111000","1111110010001111","1111110001010111","0000000100000011","1111001110111011","1111110011110010","1111101001000000","0000001101101011","1111111110101101","0000011110010110","1111100110110010","1111111111110000","1111100011100111","1111111001110010","0000000110100011","0000100110011111","1111100001001010","1111101111010011","1111110000001000","1111001010010011","1110111010110101","1111111000011010","1111100010010010","1111101011010100","0000000010110100","1111101110101010","1111101101111101","0000000010010010","1111111000110011","0000001110001111","0000000011000000","0000000110110000","1111111110011000","1111111100001001","1111111000001010","0000011000100100","0000011100010101","0000101110011000","1111100001001001","0000010101011101","0000011000001011","1111101100011100","1111100001010010","1111111101011111","1111011011100110","1111110010010110","1111100100111000","0000001110001100","1111111000111111","0000100001110101","0000001111100110","1111111100000011","0000010111000010","1111110001100000","0000000110000001","0000010100110111","1111111100101011","1111010011100001","0000000110100001","0000000110101100","0000001101110000","1111101100101111","1111111001010100","1111100100111010","0000010101100000","0000010101111110","1111110011100001","0000001110100110","1111101011111010","1111001000011101","1111011111110010","0000010111110101","0000001111011001","1111101011110101","0000011100010101","0000001111011011","1111110100110110","1111111010110011","0000001000110011","1111100000011010","1111110100011110","1111110001101111","1111110011000001","0000010011001010","0000001011111111","0000000000101100","0000010001111000","1111110101100101","1111100111010001","0000000011110000","1111101011001101","1111101011110100","0000010011101101","1111011101110111","0000001111001010","1111101100001010","1111000101011100","1111111110010101","0000010011001000","0000100100110000","1111101101100110","1111100100001111","0000001010101111","0000010101101110","0000100110000000","0000001110000100","0000011111001110","0000011101100110","0000000011011011","0000001101100110","0000000111000010","0000010010011011","0000001101011011","0000000101101000","0000011100010001","0000000101101100","0000010011000000","1111111010010000","1111100001000100","0000100011010101","0000010110000000","1111101111100100","0000001000000110","0000011011111110","1111111001000011","1111100101001010","0000000101001010","1111100110000010","0000000101100000","1111111101111100","0000001010011000","1111010011011011","1111010110111011","0000000000101111","1111101101011001","1111011101001010","1111101111100000","0000000110000100","1111101111110110","0000100010001101","0000010000111101","0000110011011010","0000000100001100","1111110011101010","0000001000000010","1111101010000100","1111110001000110","1111111010001010","0000000000011110","0000100010100110","1111010111100100","0000001011010101","0000011100011001","1111111111111011","0000011000111010","1111101010011101","0000011101100011","1111110011011000","0000011110010110","1111011000111010","1111101011010111","0001000000000111","0000001111001000","1111111110011011","1111110000010000","0000001000101010","1111011011011101","1111110001110110","1111101001100001","0000000100010111","0000000011001000","0000000000111111","0000010111100101","0000000010010011","1111111100110010","1111110001000111","0000011011011001","1111100110000001","0000100001010010","1111110011011110","0000000011001000","0000001111000011","1111110101110011","1111100111110011","0000000111000010","0000010100111000","0000011101001110","1111111111011110","0000100001011110","0000000000000011","0000001000111011","0000000000101001","1111010010001000","1111100001101101","0000011101111111","0000000010010000","0000000100100001","1111101100111000","1111111100010111","0000000110000101","1111111110101010","1111101101000111","1111110100011111","1111010000000101","0000101111110111","0000110000101001","1111000011101010","0000000100101010","1111101101101011","0000000000101111","1111110011110110","0000000011011110","1111110010010100","1111110010011001","0000100100010010","0000100100110001","0000001111010110","1111111001001101","0000100011010001","0000001000011001","0000010010100100","1111101100011001","0000011101100000","1111110011010000","0000000001101001","0000000011100101","0000000100100000","1111101011101001","0000001011000011","0000010010001100","0000000100010101","1111100010011111","1111101001111101","1111110110001110","1111101101011000","1111100100101101","0000010101011001","1111100111101011","1111101010100001","0000010111111110","0000101101101010","0000001100001000","0000110100000001","1111101101110001","0000101001111001","1111100111110101","0000001100000111","0000001110110100","0000000010000001","1111111000100110","0000100111111100","1111101100110001","0000110001111011","0000001000011001","0000100100101101","1111100101000110","0000010011000110","0000001011100111","0000000110001111","1111101100110101","1111101110010011","1111101111010000","1111100110110010","0000010111111101","1111111010100110","1111001111000100","0000011000111011","1111111001101010","0000010010111011","1111111001010100","1111110100100010","0000010110001001","1111100010001111","0000010111010111","0000100111010000","1111110101001011","1111100001010111","0000001100000000","1111100011000000","0000011101100110","1111101101111010","1111101100011111","0000010001110100","0000101110100111","0000000001100001","0000011010101101","1111111000111001","0000101001111010","1111111001010000","1111110001111110","0000110000111101","0000000101001011","0000011001001110","0000001111100100","0000010001010010","1111101100011100","0000111100101101","0000100001010110","0000001000100100","0000100110001101","1111101111101110","0000001010000001","1111111110110100","0000001100010101","1111110100111110","0000100100000011","1111101010010101","1111101101100011","1111101000000010","1111111100010110","0000000000100111","0000101100011111","1111110101110111","0000010000000101","0000000110111000","1111111111111100","1111110111010011","1111110011100000","1111101000000010","0000001101111100","0000000111101011","0000000010100111","0000010111010011","1111110111010110","0000101010010010","0000010011001001","0000011001010100","1111111101001010","1111111101111001","0000000100001011","0000100111001101","0000010111000110","0000000000110110","0000000110111110","0000010101111110","0000011100001000","0000000101111101","0000001110011101","1111110101010011","0000001011100111","1111111111110010","1111111010110110","0000011100111010","0000000000001010","0000010000011110","1111001101000011","1111111101101100","0000000101111010","0000011100010111","1111110010101001","0000011110011110","1111101011100010","1111100100110000","0000001011101100","0000010010001111","0000100010110000","1111100010000111","1111111000000110","1111100011100010","1111111000001001","0000011010100011","0000011001101010","0000000100011100","0000000001101111","0000010001111100","0000001011000100","0000001100101110","0000001100111100","0000000011011100","0000010101101101","1111110011011110","0000001011011100","0000010100100100","1111001010110100","0000010100001000","1111010101001111","1111111100111001","0000000000101011","1111101101100111","0000011100010101","0000000110110111","1111110111010101","0000010010110011","1111100111100111","0000001010101010","1111010110100001","0000001011110010","1111101001100011","0000010000100010","0000010001100011","0000000111100000","0000001111011010","0000001111101100","0000010111010111","0000000111111010","0000000001111100","1111111111000101","0000010100011010","0000001100011001","1111110011010010","0000001100011010","0000011100000111","1111110001101000","0000010111101101","0000010110101011","1111111101111010","1111101001011011","1111101011111000","0000010000000110","1111011101010100","1111110100111011","0000000001011000","1111101101101111","0000000010111110","0000001110110100","1111111100110111","0000000110001011","0000000111001111","0000100001001000","0000001110111100","0000000000000001","0000010001001110","1111111100001010","1111111100110010","0000000001010001","1111100011101111","0000000111101100","0000000100100110","0000011100001000","1111010111001110","1111111101001011","0000101010000001","0000001110100100","0000100000000010","0000000010000101","0000010111111100","0000101100100001","1111100110110100","0000011001011111","0000011010110101","1111110111101101","1111101100010111","1111101001101111","0000100110111011","1111100100001010","0000100011011100","0000100011101001","1111110000110100","1111111011110001","0000101110010110","0000001101000010","0000000011111100","0000001000000110","0000001100111001","0000000011000111","1111110010010001","1111101011010010","1111100100110100","1111010011111110","0000000111110101","0000011000011100","1111110011101101","1111101011000111","1111111000011011","0000000000001110","1111110011111100","1111111110010010","0001000010110000","0000010010010010","0000000000110100","1111110111101111","0000000001101110","1111100110110110","0000101100010011","1111100100011010","0000010000001011","0000001001000111","0000001110111000","1111101000010001","1111011100010011","1111110011101101","0000001101100111","1111110111000010","0000010100001000","1111110110111110","1111111110111001","0000011001101110","0000000110101111","1111100110110010","1111110111010110","1111101010101111","1111111011111100","1111110001100100","1111100000010000","0000001000110001","0000000011010000","0000011000111111","1111100111101001","0000001001100101","0000010011000011","0000000001110011","1111011100010101","1111101011010101","1111110110100111","1111111011100111","1111110111100011","1111110111111111","0000000000010100","0000011001011100","0000010011101011","0000001011100011","0000001010000100","0000100101011011","0000001100110111","0000001111100100","1111110110010011","0000011010110011","1111100011111010","1111011011000001","1111100001111100","0000001010111001","1111111001110010","1111111010010101","1111011101000100","1111101110111101","0000011010000110","0000001001010101","1111101110001001","0000001010101001","0000110011101101","0000110011110101","1111111111010001","1111111011011100","0000001111111101","1111100110100011","1111110101000000","1111011111111100","0000000010110001","1111110100011001","1111111111010011","0000011000111101","0000001010100011","1111111110011011","1111110101111001","0000011011000100","1111011110110011","0000100000110010","0000001100001110","0000011111110111","0000000111100010","1111101100110100","1111101111000011","1111111011101000","0000101001011010","1111010111110000","1111111000000101","1111110001000100","0000011101000111","0000010001011100","1111110100001001","1111101110000111","1111001000000100","1111100001110111","1111110001010011","1111111110011010","0000001111010011","1111100111110011","0000101011110110","0000000101011001","0000011000110001","0000111100011010","1111110101010001","1111111010101111","1111111100000011","1111110000000100","1111100101010000","1111110000110011","0000001011011001","0000000101111100","0000001010010010","1111111010111000","1111100100111010","1111111100111111","1111110000111000","1111101100101111","0000001010110001","1111110110000010","1111111001001011","0000010011110010","0000001111010100","1111100111001000","1111101000011001","1111110011111001","1111101001010011","0000000110110010","0000100101111011","0000011011011100","0000001100100111","1111101110011001","1111100110100111","0000011001110011","1111101011110001","0000000111101111","0000011100100001","1111110011100101","1111011000110010","1111011010111111","1111101110000110","0000010100000111","1111100011101111","1111011100100011","1111000110000110","0000010000111110","1111110011000011","1111111010010101","1111100100111011","1111111111000100","0000000010011110","0000000110011111","0000000011010110","1111101100100001","0000001111111000","1111111101001010","0000000001000011","1111110101110100","1111111100000011","0000001110101101","0000000110110111","1111111110111111","0000000100010011","1111110001111110","0000010010100000","1111110111101110","0000110110110000","0000000110010111","0000000100010011","1111101111100110","1111111000100100","1111111011111110","0000100001111011","1111101000111101","1111101000010000","0000001001001100","0000001011101011","1111101101001111","1111100100100000","1111110011010001","0000000010001001","0000011111001010","0000101001001111","0000000000010110","1111101110000000","0000000010001011","0000010100100100","1111100011101110","1111101100000010","0000011000001110","1111101001011011","0000001001010100","1111011000100110","0000001001001111","1111101010110001","0000011101101000","1111110010001011","1111111010000011","0000101010101100","1111110000100111","1111100010001111","0000000001101011","0000000000010110","1111011110010001","1111110011110101","0000001000111101","0000001010111110","0000000100100100","0000000111100000","0000001110001111","0000010100101111","0000000111001000","0000011110011001","1111101110110000");
	signal r_mem_img		: t_mem_img 	:= ("1111110001111101","1111111110100111","1111110110011110","1111100010011101","1111111001000101","1111100010011111","1111111110000001","0000001000111100","1111011010101100","1111110000110000","1111000010011000","1111110101010011","0000010111011110","1111101000110000","1111011010100110","0000011110000111","0000000001011101","1111111110101000","0000010001111101","1111011011001001","1111111010110101","0000000111011010","0000000101100010","1111111111001011","0000001000011101","0000010010111100","1111101111010011","0000001101011001","1111110111010000","0000000101101001","0000001010110001","0000011010011111","0000010010111111","1111101111000011","1111110110000101","0000011001001100","1111000011100110","1111101010111011","0000001110100110","0000100101101110","1111111000110010","1111101110010011","0000011101110110","0000000100101100","1111110010000100","0000010000001100","1111110100001001","0000011000011110","1111110010100001","1111111110100100","1111111011100000","0000010010110010","1111011111000011","1111011000000110","0000001010011001","0000000101001011","1111111000001001","1111100001001101","1111110110111100","0000010011111011","1111111111111110","1111101101111010","0000001111001100","0000011100000101","0000000000101110","0000010111010100","0000000010000111","0000011110001101","1111110100110000","1111111001101111","1111111111101011","1111111110101011","1111001101101101","1111111011000111","1111110010001101","1111110001001101","0000001001010101","1111110001101100","1111101101101101","1111011100100100","0000000001010011","0000010001001110","1111111111101101","1111111101110111","1111110011000100","1111111101110001","1111110111011100","1111100001111101","0000010001111111","0000000000010101","1111100100010100","1111110101101100","1111111001110000","1111111010111001","1111001101010100","0000011110110100","1111110011000000","1111011011111000","1111100101001100","1111111010100101","1111101010000111","1111111000110000","0000000000010100","1111101100110001","1111011011110111","0000000000110001","0000010011111010","1111101110110010","1111111110001100","1111111111001101","1111111010101010","1111110011110101","1111110111110101","1111100110101011","1111111001100110","0000000011000100","1111101100111010","1111110100110011","0000001001011000","0000001100110110","1111111100010100","0000001000111001","1111100000001001","0000000111010101","1111110011110000","0000000101010000","0000011001110110","1111110010000011","0000001110000111","0000100011010000","0000001000101101","1111111111111111","0000100001011100","1111111100101101","1111010110010000","0000001010001000","1111110100010011","0000001101011101","0000000011111001","0000000100000011","1111110110110100","0000001011000110","0000000100101100","0000010010001101","1111111010101010","1111011001001000","1111111111111111","0000011011111000","1111110101001010","1111110011101011","1111011011110000","1111101010011100","0000000111101111","1111100101001100","1111110000110110","1111111010110010","1111111001001010","0000010010000011","1111100000010011","0000010111110100","0000011001100000","0000001111010001","1111100011110100","0000101011001011","0000010100011111","0000001000011001","0000100010111001","0000011000110101","0000011101110110","0000100011001001","0000010101100101","0000001010101110","0000010001001011","0000011010000101","1111100110010100","1111011110001001","0000011110010110","0000011010001011","1111111000011100","0000001011101001","1111011111010100","1111101001101000","1111110101100011","1111110010110100","0000011101111001","0000100000011111","0000000100101010","0000100001101001","0000010001100100","0000011000111110","1111001100110111","1111101001110010","1111100111110010","1111010011011011","1111011000011001","0000010010010001","0000001110011010","0000000110111011","0000011010001000","1111111101110001","1111110111111000","0000011011001001","0000001110101111","0000000000110111","0000011110111100","0000001011011000","1111101011101100","1111101010000000","1111111111101001","0000000111110001","1111101010110001","0000100010100110","1111010011101001","0000001111101101","1111011001101011","0000010000101011","0000010000010111","0000011001000010","0000001011110000","0000011001101101","0000001111010100","1111110101011100","0000001010001110","1111111011101001","0000010011010110","1111111001111011","0000000101011010","0000011101100000","0000011001100100","1111110010100100","0000011011010010","0000001001101000","1111111010111111","1111110110110011","0000101000011010","0000101110001111","0000000100011101","1111101000000001","1111100111010001","1111111001100000","0000111111011110","0000001011010000","1111101010111011","1111110110001000","1111101100110111","0000000000000001","1111101010101111","0000000010111110","0000100110111110","1111011101101011","0000001111111110","1111111001110100","0000001011010011","1111101111111100","0000010100111100","0000010010111010","0000000001011010","0000001101101010","0000001010111010","1111110011111101","0000000010010101","0000000000011100","0000001101010000","1111011111001101","0000001000001010","1111101110110101","1111101101011000","1111010001111010","0000010001010110","1111110110100010","1111011111011111","0000000111001010","1111001101111001","1111110000011010","0000111101111100","1111100110011010","1111110011000110","0000011001001101","1111111111100100","0000010110110000","0000010100100101","0000010100010001","0000001011000100","1111111000111101","1111110111110000","0000000100110110","0000010000010101","0000101011101000","1111110100101011","1111011110001010","0000010100100100","0000011000100010","0000110010000010","0000100101000100","0000001100011100","0000000011111111","0000010011110000","0000001010101101","0000001110000001","1111101101001010","1111101010010010","0000001011011000","1111111010101010","1111110000111000","0000000001110110","1111101001001100","1111110100110011","1111111100111101","0000000010010111","1111010111100110","1111101010010001","1111100010100000","1111011100000101","0000000010010010","0000011100010111","1111101111000001","1111100010101101","0000010001010101","0000001101000000","0000001111100000","1111100101011010","0000001111110011","0000100001010101","0000000110011010","1111100110010000","0000001011100010","1111100010011101","1111110000011001","1111111010011001","1111110101111010","1111111011010110","1111111100001010","1111100000001011","0000011011001110","1111111100011000","0000101100011010","1111010101110001","1111101110111110","0000011111111111","1111111111100100","0000011010000100","0000001111010000","0000001010010111","1111111010111010","0000000110011111","1111011110101101","1111101000111111","0000000010111110","1111001100011100","1111110100101110","0000000011110100","1111110111000000","1111111001000100","0000000000110000","1111111101111001","1111100000101001","1111111100111011","0000000100011010","1111101101011000","0000001111001101","0000000100001000","1111010100111010","1111111111000010","1111011111111110","1111010100100010","1111111100100100","1111111010101001","0000001010111001","1111011101000011","0000000101001111","0000011011001111","1111110100110000","1111111111010010","1111101100111000","0000010000111111","1111111110100101","1111111111101001","0000000101011011","1111100110110001","1111111110110101","1111100101011011","0000000001011110","1111101001001110","0000001100111011","0000001010001011","1111011100001000","0000010111100100","1111111000001110","0000000101010011","1111111010000101","1111000010101101","1111010111101101","0000000011101001","1111110110001101","0000011111110011","1111111110000110","1111101110101011","0000000111011011","1111111011110111","1111110010101001","1111111101010101","0000010000110110","0000001111100000","0000000110011010","1111110011000100","0000001110100000","1111111101110101","0000000001001110","0000011111000001","1111110000001101","1111110011110110","1111111000100011","0000000101101111","0000000000110111","1111010101111010","1111111001111000","1111101110010111","0000010000110101","1111110010010001","0000100111001100","1111101101110110","0000101110111001","0000001001101011","0000000110111010","0000001011001011","1111111000010000","1111111110100011","0000001011101110","0000001011101100","0000001101001110","0000010101101111","1111111111110101","0000001001000001","1111100101000110","0000000101100001","1111100101001110","1111101001111100","1111111100010111","0000000111101001","1111101101110011","1111101001011111","1111110110000110","1111111111011011","1111111111110011","1111111001000000","0000000000000000","0000001110101101","1111110110100011","1111111100000011","1111101001010001","0000010001000110","1111110101011001","0000011100001011","0000010010011001","0000010111001011","0000011000001111","0000001010100100","0000001010110110","0000010010100010","0000001010101000","1111011001011001","1111010111101100","1111101001101100","0000000100011111","1111011011010111","1111110100011111","1111101000101000","1111110011000010","0000101000011010","0000000100110010","1111110010111000","1111101111100011","1111111001101010","1111100010001101","0000011100100110","1111110100010111","1111100101100100","1111110110111011","0000010011101110","0000000110110101","1111111101001000","0000000010111000","1111101111000000","0000000000000000","1111101011010001","1111110010111111","0000000001100110","0000000111000100","1111100011010111","1111011000011110","1111100110010110","0000010010011010","0000011010110001","1111110010110101","0000001011001100","1111111101110001","1111110110001001","1111110111010110","0000000011111101","0000001001111100","0000011000101101","1111110100110111","0000011100110001","0000000101011010","1111111101000010","0000000101101101","0000010001110010","1111110010010101","0000100101110001","0000010000001010","0000000010101010","0000000011011110","1111111000111000","1111101111100000","1111100011000111","0000011011100011","1111110011000001","1111100100001001","1111100010000111","1111111100111111","1111110011010011","0000010011001110","1111101101101100","1111110101011000","1111011111110011","1111100110100110","1111101111010000","1111101100000101","1111000010011000","1111100110110110","0000000110011110","1111100101011111","0000000100101101","1111101000011000","1111011111001010","1111100110110110","0000000110111011","0000011101010101","1111111011101111","0000001000110110","0000110000100001","0000010001000011","0000011111101011","0000001001010011","0000001111111000","1111010101011100","1111111101011000","0000001011100010","0000000011010110","1111111110010001","0000010110100011","0001000100100001","1111101110111101","0000011100011111","0000000110101110","0000000101111101","0000010000001100","0000001100001111","1111011110101010","0000011010111011","0000010011110001","1111111100111011","0000010011111011","0000010000010001","1111110101010010","1111110010000001","0000000000100010","0000010101011101","1111011101101001","0000001100000000","1111011111101011","0000001001100000","1111111011100100","0000000100000001","1111100001000011","0000100001110000","0000011000011101","0000001010000000","0000010001100101","1111110100111110","0000001100010111","0000010101100011","0000001111111111","1111110111000111","1111111011110010","1111111110001010","0000101000001011","0000100011111001","0000011001000011","0000100000011111","1111101101111100","0000010011111101","0000000000111111","1111110111101111","0000011111111010","1111100111110001","0000011100100011","1111110100110101","1111101111101110","1111111010110110","0000001100011000","1111101001111111","1111111101001011","0000001010111001","1111100011000111","1111010101000111","0000000011010010","0000011010011000","1111111100011010","0000011110110100","1111011001100011","0000000000000010","0000000101110010","0000000010011010","1111110111100010","1111110101001111","0000000100001110","0000011100010010","0000010101110110","0000001001000010","1111100111001011","0000001011010011","0000010100100110","0000100100000101","0000001011000011","1111101001001000","0000011111100010","0000001100000010","0000011110101000","0000000111100000","1111110111011100","0000010000100111","0000011111110110","1111111110101010","1111111001100010","1111110111011000","0000010111100110","0000000010010101","0000001101010000","1111101001011111","1111110000111011","1111110000010000","1111110110101001","1111111101011110","0000001111101001","0000100110100010","1111110111110001","0000100011101110","0000001100111011","0000000011110010","0000011000101101","0000100101011110","1111111000000000","0000001010011111","0000001101101010","0000101010111111","0000011001010011","0000011001000100","0000101110001011","1111110010011010","0000001001011000","0000010111110011","0000000000111110","1111110000000011","0000011101110011","1111100001010100","0000011001000101","1111110010000111","1111011001000101","0000001011101010","1111111100010011","1111111100011001","0000001101101100","1111011111001110","1111110100001101","0000011010110001","1111111000101011","1111100001000100","0000000011010100","0000001110010111","0000011000100010","0000000110111101","1111110011111101","0000011100001010","1111100011110100","1111111001010001","1111110101111001","0000001010001001","0000001111010100","1111111101111001","1111100010000110","1111100101011011","1111101100100011","0000011001101110","1111101000011000","1111111101000100","1111100001001010","1111110110001111","1111111101001001","1111111110010111","1111111100100001","1111011101010000","1111111001011100","0000000101001101","0000011001011001","0000010101000000","1111111011110101","1111111010000111","1111110011110001","0000001001100000","0000001111100111","1111100111111010","1111111110001000","0000000000110101","0000011111110111","1111111110010100","1111110010000000","1111111011111000","1111111001001100","0000000100000000","1111111011010111","0000101110110001","1111011110110001","1111101111010010","0000011000111011","1111111101100001","1111101111001001","1111111010011111","0000010011010110","0000110011110101","1111110010011000","1111011011011100","0000100100101011","0000010010001111","1111011100011010","1111010110111000","0000000101110101","1111111111010000","1111101111101000","0000000110000001","1111100101101101","1111101111101010","0000001111111010","1111110011110000","0000010111111000","0000000000001010","1111111111110110","1111111101010100","1111111001110001","0000011110000010","0000100111011001","0000001010111111","0000011100110010","1111011011010111","0000000111001110","0000000110110000","0000001000100110","1111111101110101","1111100010101100","0000000101000000","1111111000100011","0000011001001110","1111010010111011","0000010111011010","0000000010111100","1111001101100100","0000000011100111","1111101001111101","0000110011111101","1111111011111101","0000001110011101","1111110110011110","1111111010111100","1111110000010000","1111110101111101","1111111100101101","0000101010000100","1111100111001111","1111100110000111","0000000110010100","1111010110110010","1111101111001011","0000001001101001","1111110101001001","1111110110101110","1111110100011110","1111011000100011","0000000001011100","1111100111101101","1111111000010101","1111110001001100","0000001100001110","0000100000000110","1111111100101100","1111101010111011","1111101101011010","1111111110101111","1111101010010001","1111101111010111","0000001111001100","0000000111111101","1111101111001001","1111111100000000","0000010000011110","1111110001101101","0000000110100100","1111100110110101","1111110001110001","1111010100111101","1111011001111011","1111110010100000","1111101001000011","1111101001100001","1111011001100010","1111101110111001","0000001100010110","1111100011100100","0000101010001010","0000001011111110","1111011101111100","1111111101110000","0000001000001001","0000000100010001","1111101011111001","0000001110100111","0000000001111010","1111110101011010","1111110100100100","1111111101110000","1111001111010111","1111100111000101","0000001000000000","0000001010100101","0000000101000100","1111110000111110","1111111010010110","0000011011101111","0000101110001111","0000000000111000","1111111110110001","0000001011110111","0000001010110111","0000000110111011","1111111100100100","1111101010101001","0000010100101111","0000100000110111","1111110101000010","1111001100111101","1111110110000100","1111110010100010","1111101110010001","0000001101011000","0000001011110010","1111101001110101","1111111001100101","1111100101110000","1111100000110010","0000000011110111","0000001110111011","0000000010000111","1111110100010001","0000010101110011","0000001010010000","0000001111001010","0000001100001001","1111111100100111","0000001110010110","1111100000100001","1111110100100111","1111111011011101","1111000110001110","0000000010110000","1111110001101110","1111101001110011","1111111010000011","0000000111111000","0000010110000010","0000011100011100","0000011000011000","1111110110100011","0000100010011110","1111011000111111","0000100010101001","0000001011000010","0000000101111110","0000001100111011","0000000100101010","1111110010001010","0000010011111001","1111101010110100","0000100011011110","1111111110011010","0000010110111100","1111100110000111","1111110010110111","0000000010011100","1111111100111100","1111101100111001","1111010111010110","1111111001111001","1111110011111010","0000010100001000","1111100011101100","1111111101010101","1111111100100100","1111111101001001","1111111001101000","0000010000101010","1111000101111110","0000001100110000","0000001000100110","0000000101101010","0000111100110000","1111100111100000","1111110101110100","1111111110011010","1111100000000100","1111111001001001","0000001101011101","1111111100001110","1111111011101110","0000011101011000","0000000010010101","0000110100001110","0000000100011000","0000001100100000","0000001000111101","1111110011111000","1111111001100101","1111101010011011","0000010010011000","0000110111111011","0000010001010110","1111101011010110","0000001011001000","0000011110000011","0000010110111000","1111111000010000","0000011010011101","0000011010100101","0000001001010011","0000000010010110","1111100111111110","1111011111110100","1111110010011101","1111100110110001","1111111000010101","1111101011001001","0000010111101110","1111111001000010","0000101111101010","0000100101010001","0000010100100101","0000001000100100","0000000110011011","1111101010011110","1111110001001000","1111110000001110","1111100110111110","1111101011111100","0000000101101010","1111101000001000","1111111111001010","0000010110011111","0000100111010101","1111100101110011","0000000111101110","1111111100011011","0000000100100110","1111011101001010","0000100101100110","0000101010001101","1111110111101000","0000100100111011","0000011100110001","0000101110101000","0000001100000101","0000001110011001","1111110001010110","0000011011110000","0000100110111100","1111100011100101","0000011100111111","0000100111110110","0000010111110000","0000011001101010","0000011110110010","0000010000000100","0000110001010100","1111111010101000","0000000011001111","0000010101101111","0000001010010011","0000010101111001","1111011011110011","0000001000110011","0000110001110000","0000001000100010","1111011011110100","0000000100010010","0000001100001000","1111101100011100","1111110110011111","1111110011100001","1111100111101000","1111111110001111","0000000110001101","0000011010000010","1111110001101110","0000010010111001","0000011010110111","1111101010000001","1111110110011011","1111110010001000","1111100111111000","1111101010100101","0000000100011100","1111110101101100","1111101011010100","1111011000011101","0000010010011111","1111101111011010","1111100010100001","1111100110111110","1111101011010111","1111111101100000","1111001001010010","1111110100011010","0000010001000111","1111101100001111","1111101001000001","1111100111001101","0000111010111001","0000000010000110","1111110010110110","0000001000101000","0000000001100001","0000010111011010","0000011011101010","0000100000000001","0000010001010110","1111111010001100","0000001111100011","1111110010000100","0000001110100100","1111111001000110","0000100011000001","0000001010010001","0000001101111101","1111111011101000","0000101000110101","0000010001101011","0000001011011001","0000110100010001","0000100100111101","0000001101111010","0000000010000101","0000100100110100","0000001010101111","0000010010101110","0000100010101100","0000100010100111","1111111001100000","1111111100010010","1111110100010100","1111010001100110","0000000110011010","0000001010001100","1111111110001000","0000000010001001","1111110101111011","0000010110100111","0000001100001111","1111010011101010","1111101100010000","0000001101000011","1111110101110111","0000011011100111","0000010111011000","0000001101100010","0000000001111011","0000010000100010","0000000010101001","0000001001001111","0000001010100010","1111110010100001","0000001111011101","1111111000001111","0000000000100011","0000001000010010","1111111000001101","0000001011000010","1111111000100001","0000101101110101","0000011001001010","0000110001110001","1111111101100001","1111111001110111","1111110101000110","1111111110000011","0000000111101000","1111001000001011","1111111000011001","1111110001101100","1111101101110100","1111100111100101","1111010101111000","1111101111000001","1111101010110011","1111010011011110","1111101001101101","0000001100101101","1111011000001000","0000000110100000","0000010001111100","0000000101010000","1111100001000000","0000010001100110","0000001111111101","1111111011001111","0000000111100100","0000101110001001","0000100000101101","1111110011000010","1111110111000111","0000010110101011","1111100110000001","1111110110110000","0000010011011111","1111111101001101","0000001000011100","0000010010101011","0000101010110111","0000000101000110","0000110111011100","0000001100011101","0000010011010001","0000110000001101","0000001101010111","1111110011110011","1111111011111000","1111111101101100","1111110010011010","0000001011111111","1111010111011011","1111101101110010","1111101010011101","0000000110110010","0000000000000100","0000000010110001","1111111101001101","0000001001100101","0000010010110111","0000010011110010","0000001100010000","1111111011000011","0000010000100111","1111101110100110","0000001000010110","1111111011000111","0000010111010110","0000001001001000","0000101100010001","1111100010100101","1111001011100011","0000001110101011","1111111001101100","0000000111100001","1111110011101110","0000000001110111","1111111101011010","0000000011101100","0000000001110111","1111111111101000","0000010010001001","0000010101010011","0000000010110000","0000010000100000","0000000101111001","0000101000010110","0000000100101110","0000110001100000","0000001011110101","1111100101010111","1111100001110110","1111010010011100","0000100000010011","0000011101101110","0000001000111100","1111010011000110","0000001111110101","1111100110101101","1111011011111100","1111100010100101","1111011011000000","0000011010100110","1111100011101010","1111011101111110","1111111100001000","1111101111100111","1111111010011100","1111111010001000","1111110111000110","0000011001100001","0000101110110111","1111111101011101","0000000001101100","0000000011101101","0000001001011001","0000000010001000","0000110011101111","0000000101000100","1110111110000110","0000010110101011","0000000110100111","1111100011001111","1111111101100101","1111111101011010","1111100010111101","1111110110001111","0000010110000110","0000000001101110","0000001010100011","1111011101111100","1111010011000110","1111010011100100","0000010000110101","1111100100000000","1111111000110001","1111111111100001","0000010010001100","1111101100100100","0000010101011010","1111110010100000","1111111100111100","0000001100101111","0000010110011010","0000011101011101","1111001001100010","1111111110011110","1111111001100000","1111110000011000","0000010011001000","1111110001010111","1111101101101000","1111110011000110","0000000001111010","1111111001101101","0001000000100100","0000001100100100","0000101010111110","1111110010000011","1111101110101111","1111111110111000","0000000101000010","1111101010110101","1110111101001110","1111101000001111","1111101110111101","0000001101110111","1111110010111000","0000010110001010","0000000110101110","0000001000100100","0000001000011011","1111110101001101","0000001001110100","0000110000101010","0000100111011111","1111110011110111","0000000000111000","0000011000101111","1111110100011001","1111110110011010","1111111110100001","0000010100011000","1111110110111000","0000001001001100","1111110010110001","0000100100010100","0000010001011000","0000110010111000","1111111000101110","1111111100000010","0000010110110010","1111110110000100","0000111001010010","1111111111011101","1111101011101011","1111111010001000","0000110101101011","0000010110100110","0000010110000000","0000101011010000","1111111111101100","0000001000001111","1111111011110011","1111111110110101","0000011101000011","1111111111011001","1111111010011010","1111110100010101","1111101111101011","1111011000010100","1111000101010110","1111100100001000","1111101111100100","1111110110110101","1111101110010110","0000000110110111","1111110011011001","1111111001101110","1111110011000111","1111011101101110","0000011010110111","1111011111100011","1111100101110111","1111111011111110","0000100100000111","1111110000001101","0000000110000000","1111111011001111","1111100010110001","0000001100110111","1111111111101001","0000001010011100","0000001100011010","0000000101001111","0000010001001110","1111111011111110","1111110011101010","1111101111100111","1111101100101111","1111101111101000","1111111001001000","0000000000010000","0000001000110011","1111100110101110","1111111110011010","1111111011011010","1111101100111110","1111101110101111","1111111010101001","0000011000111110","1111111010001111","0000001110010100","0000110011000000","1111100011011100","0000010101110011","0000011111010101","0000011000111101","0000011001100011","1111110101100000","1111100101000101","1111101001100001","0000000101110100","1111110100001101","1111110011111001","1111101000000000","1111010111101001","0000100011111101","1111101100010110","1111100000001000","1111110001110001","1111111010000100","0000100101100100","0000011110100110","0000011101100100","0000100110100011","1111111000101011","0000001111000001","0000000111001101","0000000101100110","0000010011001100","0000010110000101","1111110110100001","0000001011000000","0000010110100100","1111111001101011","1111110101000000","1111011111101101","0000100011110001","1111110000011111","1111111011011100","0000010110010111","1111110010010111","1111101110110000","0000000111001100","1111100001101101","1111001000001110","1111111101000110","1111111101111100","1111011010010110","1111001000000000","0000010000111111","1111110010110111","0000000111011001","0000000100010101","0000100010110011","0000010000000110","0000000111010001","1111111000010000","0000001010000000","0000011110100010","1111001111111101","0000000010000100","1111001111010100","0000001010010100","0000000011011100","0000001001010110","0000001011111100","1111011101011010","0000010000000100","1111101111101100","0000011100111010","1111111100110100","1111100110111011","0000100111111011","0000010011110110","1111110111110001","0000010000000010","0000001000001110","1111111011011010","1111100000001101","1111110000111101","0000001110100100","0000000000111101","0000001110100011","1111110110011111","0000011001100110","0000010011110000","1111111111011100","1111101011100111","1111100001101000","0000000010001111","0000010010110001","1111111101011110","0000010010111000","1111100110000110","0000010010110001","1111110001101101","0000000001100101","0000001010101101","1111101100110010","0000000100000110","1111010110000011","1111110000011000","0000000010100001","0000100010000011","0000011010001111","0000000100010100","1111111011100111","0000101100111000","0000100101011111","0000100010111101","0000001000100011","0000101001111010","1111110111001000","1111110001011010","1111111110010101","1111110001100000","0000001100010110","0000000011011011","0000001101111011","0000000100011001","0000000111100001","0000010111011001","1111100100110100","0000101110111000","1111111110100000","1111111111001011","0000011100111010","1111111111111110","0000011000011100","0000110110111111","0000000101001000","1111110101110010","1111100110001000","0000100000010001","0000110100100101","0000101010001011","1111111001101101","1111100000001001","1111101111100110","0000011010000110","0000000001000101","0000010011000111","0000000100100011","0000010101000000","1111100111101011","0000010110100001","1111111011000111","0000000101110011","1111010111101011","0000100101110100","1111100111010011","1111101000011111","0000001000011000","0000000000111001","1111011111010001","0000001100101001","1111100110101101","0000000001011111","0000001000111000","0000010011100000","0000000111111111","1111111100101010","1111100100111101","1111011101101110","0000001001100101","1111110111001000","1111110111111100","1111111010011100","0000000000011101","1111100100111111","0000000011010101","0000001110110110","1111010111101010","1111111111110011","0000100101111011","1111110101010101","1111100100110111","0000010001000111","0000000111001100","1111110111110100","1111110111011111","0000010100111001","1111101001110101","0000000101001110","1111101100111001","0000000110011110","0000010110001110","1111011011100001","1111100111100111","1111111000101100","1111011111100100","0000100011010110","0000010011100001","0000000010010111","1111111010101001","1111100010100100","0000000001110111","1111110111010110","1111100001101011","0000010100011001","0000000010001100","1111101101111111","1111111001100010","0000001000111000","0000110101011001","0000010100001010","0000010011110011","1111101100111101","0000000111110111","0000011101011010","0000000111101110","1111101111100000","0000000100010000","0000010110011111","1111100011100000","1111111110100101","1111110101001100","1111100001001010","1111100100110110","0000001111111110","0000101011111110","1111100111101001","1111111001011001","0000001111111001","1111101010100110","1111110010000000","1111110110110100","1111101110011011","1111111100001101","0000011011101001","1111110111001100","1111010011001011","1111111101110101","1111010000100011","1111011000010101","1111101111100011","0000011000010001","1111100000010110","0000011011110110","1111011101011000","0000011100011001","0000000100001001","1111110010000001","0000001100110001","1111110100010111","0000000110101111","1111110000110100","1111100011001101","1111011010001011","1111110100101111","0000000101010011","0000000100011001","0000100010011001","0000011001101111","0000011101110010","0000101010011011","0000011100001101","0000011011000000","1111101111101011","0000001101001000","0000100001011100","0000000111000000","0000000111011110","0000000000111110","0000001000000000","0000000010100011","0000000010011001","0000000110101000","1111101100011001","1111101010100011","1111101001000111","1111100100011000","1111010100101110","0000100100001001","1111110001001011","0000000000100110","1111111100010001","0000001011000010","0000100001000111","0000011111101001","0000010011000010","1111101101100011","0000100100001100","0000000000010010","1111101011111110","0000000100010100","1111010101000000","1111100101110010","1111100101011110","0000001000101100","1111110100000001","0000011101000111","0000100101101001","0000011011111001","1111101010001011","1111001001100100","1111101111010001","1111100010101100","1111111011010111","0000010001110101","0000010011000110","1111111010110000","1111111011000100","1111101000011101","0000001010000000","0000010110110011","1111011101101000","1111110011000110","0000000111001100","0000001010001010","1111101110010011","0000100010100110","1111111000010110","1111111101100100","0000000010111110","0000000101101000","1111010101011001","0000010100010011","1111100001000101","1111010001011000","0000100000000010","1111011000001100","1111111110110111","0000001001110110","0000100011010110","0000011010101100","0000101100000010","0000001001011100","1111111111101000","0000001101000010","1111110110000000","1111101101111110","1111101010101011","1111100101110111","0000011101001000","0000010101101110","1111100100101010","0000011100001010","1111111001010011","0000000101101101","1111101000000100","0000000011110101","0000100100100010","0000011010000010","1111101111100100","1111111111001011","1111110001111000","0000001111011011","1111111100101100","0000001001010011","0000010101101000","1111111001000110","1111110101010011","1111110111110001","0000010101001101","1111101110111011","1111010100011111","1111010111101001","1111011101111100","0000010010010001","1111101111111100","0000001110101110","0000001011111110","1111010100101010","1111010100100111","1111110110001001","1111111111010110","1111100100111101","1111110101100001","0000110101000101","0000000010110001","1111111101000111","0000011001001011","0000001001010001","0000001110001111","1111011101100111","1111111101011100","1111111011100101","1111111111010010","0000000000000110","0000000000111010","0000011110101100","0000111001110101","1111110011001110","0000100001000000","0000000101110110","0000001111100111","0000011011101100","0000000010111010","1111010110000101","0000011001010011","0000010111110011","0000000110101101","1111101011101010","0000101101011000","1111110111011000","0000001011000101","0000000011110010","1111011001100110","1111100110111110","0000000110011001","0000010011101000","0000011101011110","0000000001000100","0000001101111010","0000101010001010","0000000101100101","1111101101110100","0000010101001001","0000011100001011","1111101101001110","0000000001100010","0000001001111101","0000011000001110","1111111000010001","0000010011101011","0000010000101010","0000010011100101","0000011100111100","0000010110100001","0000110100100111","0000001100010001","0000001110101110","0000101010000001","0000100110011001","1111110011110010","0000001111100011","0000100001001101","0000000000010101","1111111000111010","0000000001100000","0000010100000000","1111101001010001","0000010111011010","1111110110001111","0000011000111110","0000000001011010","0000010011000110","0000001011010110","0000000001011001","1111101101000010","1111110111000111","1111100101110111","0000010110100111","1111011010110101","1111111100110001","1111101001111011","1111100011101101","0000001011111111","1111101000111000","1111011111001110","1111101001110110","0000010111001101","0000001111001111","0000100011101110","1111111100001111","0000000011010011","0000100110000100","1111111010111000","1111110010010110","1111110000011100","0000101011110001","0000101010101111","1111111011000001","1111111010010110","0000000100111001","1111101011110001","0000010100010011","0000001101011011","1111101001101000","0000000111100111","1111110011001101","1111110100110010","1111000100011100","1111100111111011","0000011100110110","0000100001011111","0000101100110001","0000001000101001","0000010001010011","0000000000011001","1111101101101011","0000001001111100","0000001101000100","1111010101111100","1111110110011100","1111111011001110","0000001010000110","1111111110111001","1111001001001001","1111111001010101","1111100101011000","0000001010010101","1111101111111101","1111010101111110","1111100110101100","0000111001100001","0000000000110110","1111111010100110","1111110101010101","0000001110101100","1111111000110000","1111010101000010","1111111111010100","0000100010000010","0000001000001101","1111110011110000","1111011101100010","1111101011110001","1111111001100101","0000011001100011","0000001101010000","1111110100111001","0000001010111100","1111110001001001","1111111001101111","1111101100011110","1111110111010011","0000010010011001","1111111010010010","0000010010101000","1111000001100110","0000100110111101","1111011001111110","0000001100100100","1111110000111111","1111000110111110","1111100100010011","0000011001011011","1111111100110000","1111100101010011","1111101000000010","0000100000101110","0000000010110111","0000010011011101","0000100110000000","0000001111000010","0000100110000101","0000010010010011","0000001111001100","0000011001100100","1111100100000000","1111101010111100","0000010100011100","0000011111000000","0000010001111010","0000011001010110","0000100001101110","0000001101101110","0000101010111001","0000010110100100","0000001110011011","1111001111010100","1111010011111110","1111010100110000","0000000011101000","0000001000111101","1111101000000001","1111101111100011","1111011100011000","1111100010000100","0000000001000000","1111011100000001","0000110001100000","1111011011100010","1111111010110101","0000011100110101","0000001101110011","1111111111100100","1111111011010010","0000000111100111","1111111110010100","0000000000010111","1111010011011001","0000000000111111","1111011100010000","1111111010011101","1111001101100111","1111111110111101","0000000001000001","1111110110110011","1111101110011100","0000000000010011","0000101110010010","1111101100100101","0000001101110110","1111110000100111","0000100110110000","1111111000001001","0000000010110111","1111110011001001","1111111110110111","0000100100110110","1111111101010111","1111010110100100","1111111101000101","1111110100100011","1111101111000001","0000110010101000","0000000111011100","0000001100111110","0000000101100100","1111101110101010","1111111001110010","1111111000100111","0000000010101111","1111100111100000","0000001101010000","0000000000101001","0000011100011100","0000000101100100","1111110101010110","1111111011100110","1111010101111011","0000010011111100","0000100010001000","0000000011001110","0000000000001100","1111101110010010","0000000101000100","0000000110111101","0000011001101110","1111111110101000","1111110011010111","1111110111111011","0000001111010000","0000001011011111","1111110100010011","1111100100000101","1111110011000011","1111111111100110","1111111001011000","1111011111101001","1111100010001100","0000000111110111","1111111110100011","0000100001110011","0000010001010100","0000110000010110","0000000100001000","1111110000101011","0000001000011001","1111111000111111","0000011110010100","1111100011010010","0000001000011001","0000001011101011","0000000010100001","0000000000100010","1111111101001110","1111101110110110","0000000100010100","0000000001000101","1111110100001100","0000011001001010","0000011101010111","0000000010001110","0000010101000110","0000101101010100","1111011101110110","1111111000100100","1111110100011010","1111111000110000","0000001000100000","1111110110000110","1111110101100001","0000001010000100","0000000011010100","0000001001111011","1111110011110110","1111100001000101","1111110011110000","1111101100110000","1111110000101011","1111011000110000","1111101100111000","0000011111010110","0000001111111011","1111101101000011","0000010011001101","1111111011111110","0000110001110011","1111111111010101","1111101110000000","0000001100111100","0000010001100111","0000011001100101","1111101001011110","0000011010111110","1111111010100010","0000000100111001","1111110000110100","0000000010110111","0000000100001110","1111111110111101","0000001010001000","0000100000100010","1111111110010100","0000000101011100","1111101110010000","0000011100110100","0000010100011010");
	signal r_mem_abs		: t_mem_abs	 	:= (others => (others => '0'));
	signal r_mem_cn_abs 	: t_mem_cn_abs := (others => (others => '0'));
	
	-- ABS signals
	type t_abs_sm is (s_idle, s_process, s_write, s_done);
	signal r_abs_sm		: t_abs_sm 	:= s_idle;
	signal r_abs_enable	: std_logic := '0';
	signal r_abs_index	: natural range 0 to g_frame_size := 0;
	signal r_abs_done		: std_logic := '0';
	signal r_abs_done_all: std_logic := '0';
	signal r_abs_real 	: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_abs_img	 	: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_abs_result 	: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	
	component abs_complex is
		generic(
			g_bits			: natural := c_bits;
			g_fxp_high		: natural := c_fxp_high;
			g_fxp_low		: integer := c_fxp_low);
		port(
			i_clk				: in std_logic;
			i_enable			: in std_logic;
			i_real			: in std_logic_vector(g_bits-1 downto 0);
			i_img				: in std_logic_vector(g_bits-1 downto 0);
			o_done			: out std_logic;
			o_complex		: out std_logic_vector(g_bits-1 downto 0));
	end component;
	
	-- Mean signals
	type t_mean_sm	is (s_idle, s_process, s_done);
	signal r_mean_sm			: t_mean_sm := s_idle;
	signal r_mean_enable		: std_logic := '0';
	signal r_mean_rst			: std_logic := '0';
	signal r_mean_input		: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_mean_result		: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_mean_index		: natural range 0 to g_frame_size := 0;
	signal r_mean_done		: std_logic := '0';
	signal r_mean_done_all	: std_logic := '0';
	
	component mean is
		generic(
			g_bits			: natural := c_bits;
			g_fxp_high		: natural := c_fxp_high;
			g_fxp_low		: integer := c_fxp_low;
			g_frame_size	: natural := c_frame_size);
		
		port(
			i_clk		: in std_logic;
			i_enable	: in std_logic;
			i_rst		: in std_logic;
			i_input	: in std_logic_vector(g_bits-1 downto 0);
			o_result	: out std_logic_vector(g_bits-1 downto 0);
			o_done	: out std_logic);
	end component;
	
	-- Standard Deviation of the Centered Normalized Instantaneous Amplitude signals
	type t_std_cn_sm is (s_idle, s_divide, s_read_abs, s_abs, s_std, s_done);
	signal r_std_cn_sm 			: t_std_cn_sm := s_idle;
	signal r_std_cn_rst			: std_logic := '0';
	signal r_std_cn_enable		: std_logic := '0';
	signal r_std_cn_input		: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_std_cn_mean			: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_std_cn_pdone		: std_logic := '0';
	signal r_std_cn_result  	: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	signal r_std_cn_done			: std_logic := '0';
	signal r_std_cn_done_all	: std_logic := '0';
	signal r_std_cn_index		: natural range 0 to g_frame_size := 0;
	signal r_cn_abs				: sfixed(g_fxp_high downto g_fxp_low) := (others => '0');
	signal r_temp_cb_abs			: std_logic_vector(g_bits-1 downto 0) := (others => '0');
	
	component standard_deviation is
		generic(
			g_bits			: natural := c_bits;
			g_fxp_high		: natural := c_fxp_high;
			g_fxp_low		: integer := c_fxp_low;
			g_frame_size	: natural := c_frame_size);
		port(
			i_clk		: in std_logic;
			i_rst		: in std_logic;
			i_enable	: in std_logic;
			i_input	: in std_logic_vector(g_bits-1 downto 0);
			i_mean	: in std_logic_vector(g_bits-1 downto 0);
			o_pdone	: out std_logic;
			o_result	: out std_logic_vector(g_bits-1 downto 0);
			o_done	: out std_logic);
	end component;

 begin
	
	complex_abs_compoennt	: abs_complex port map(i_clk, r_abs_enable, r_abs_real, r_abs_img, r_abs_done, r_abs_result);
	mean_component				: mean port map(i_clk, r_mean_enable, r_mean_rst, r_mean_input, r_mean_result, r_mean_done);
	std_component				: standard_deviation port map(i_clk, r_std_cn_rst, r_std_cn_enable, r_std_cn_input, r_std_cn_mean, r_std_cn_pdone, r_std_cn_result, r_std_cn_done);
	
	p_complex_abs : process(i_clk, i_enable)
	begin
		if rising_edge(i_clk) then
			case r_abs_sm is
				when s_idle =>
					r_abs_done_all <= '0';
					if i_enable = '1' then
						r_abs_enable <= '1';
						r_abs_sm <= s_process;
					else
						r_abs_sm <= s_idle;
					end if;
				
				when s_process =>
					if r_abs_index < g_frame_size then
						if r_abs_done = '1' then
							r_abs_sm <= s_write;
						else
							r_abs_real 	<= r_mem_real(r_abs_index);
							r_abs_img	<= r_mem_img(r_abs_index);
							r_abs_sm		<= s_process;
						end if;
					else
						r_abs_sm 		<= s_done;
					end if;
					
				when s_write =>
					r_mem_abs(r_abs_index) <= r_abs_result;
					r_abs_index	<= r_abs_index + 1;
					r_abs_sm		<= s_process;
				
				when s_done =>
					r_ft_state(0)<='1';
					r_abs_index    <= 0;
					r_abs_done_all <= '1';
					r_abs_enable <= '0';
					r_abs_sm			<= s_idle;
				
				when others => 
					r_abs_sm <= s_idle;
					
			end case;
		end if;
	end process p_complex_abs;
	
	
	p_mean : process(i_clk, r_mean_enable)
	begin
		if rising_edge(i_clk) then
			case r_mean_sm is
				when s_idle =>
					r_mean_done_all <= '0';
					if r_mean_enable = '1' then
						r_mean_sm <= s_process;
					else
						r_mean_sm <= s_idle;
					end if;
					
				when s_process =>
					if r_mean_index < g_frame_size then
						r_mean_input <= r_mem_abs(r_mean_index);
						r_mean_index <= r_mean_index + 1;
						r_mean_sm	 <= s_process;
					else
						r_mean_sm <= s_done;
					end if;
					
				when s_done =>
					r_ft_state(1)<='1';
					r_mean_done_all <= '1';
					r_mean_sm 	<= s_idle;
					
				when others =>
					r_mean_sm <= s_idle;
					
			end case;
		end if;
	end process p_mean;
	

	-- Standard Deviation of the Centered Normalized Instantaneous Amplitude
	p_std_cn_inst_amp : process(i_clk, r_ft_state)
	begin
		if rising_edge(i_clk) then			
			case r_std_cn_sm is
				when s_idle =>
					r_std_cn_done_all	<= '0';
					if r_ft_state(1 downto 0) = "11" then
						r_std_cn_enable <= '1';
						r_std_cn_sm <= s_divide;
					else
						r_std_cn_sm <= s_idle;
					end if;
				
				when s_divide =>
					r_std_cn_enable <= '0';
					if r_std_cn_index < g_frame_size then
						r_mem_cn_abs(r_std_cn_index) <= to_slv(resize(to_sfixed(r_mem_abs(r_std_cn_index), g_fxp_high, g_fxp_low) / (to_sfixed(r_mean_result, g_fxp_high, g_fxp_low)-1), g_fxp_high, g_fxp_low));
						r_std_cn_sm		<= s_read_abs;
					else
						r_std_cn_index <= 0;
						r_std_cn_sm	<= s_std;
					end if;
					
				when s_read_abs =>
					-- Why is it necessary to use the quotes in abs function?
					r_temp_cb_abs 	<= to_slv(resize("abs"(to_sfixed(r_mem_cn_abs(r_std_cn_index), g_fxp_high, g_fxp_low)), g_fxp_high, g_fxp_low));
					r_std_cn_sm		<= s_abs;
				
				when s_abs =>					
					r_mem_cn_abs(r_std_cn_index) <= r_temp_cb_abs;
					r_std_cn_index <= r_std_cn_index + 1;
					r_std_cn_sm <= s_divide;
					
				when s_std => 
					r_std_cn_mean <= r_mean_result;
					if r_std_cn_index < g_frame_size then
						if r_std_cn_pdone = '1' then
							r_std_cn_input <= r_mem_cn_abs(r_std_cn_index);
							r_std_cn_index <= r_std_cn_index + 1;
							r_std_cn_sm		<= s_std;
						end if;
					else
						r_std_cn_sm <= s_done;
					end if;
					
				when s_done =>
					r_ft_state(2)<='1';
					r_std_cn_done_all	<= '1';
					r_std_cn_index 	<= 0;
					
				when others =>
					r_std_cn_sm <= s_idle;
					
			end case;
		end if;
	end process p_std_cn_inst_amp;
	
	r_mean_enable <= r_abs_done_all;
	o_done <= r_std_cn_done_all;
	
	o_ft_0 <= (others => '1');
	o_ft_1 <= (others => '1');
	o_ft_2 <= r_std_cn_result;
	o_ft_3 <= (others => '1');
	o_ft_4 <= (others => '1');
	o_ft_5 <= (others => '1');
	
 end bhv;