library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library amc_library;
use amc_library.data_types_pkg.all;

entity ram_l2_n7 is
	generic(
		g_width   : natural := c_bits;
		g_depth 	: natural := 50;
		g_addr_bits : natural := 5);
	port(
		i_clk			: in std_logic;
		i_wr			: in std_logic;
		i_addr		: in std_logic_vector(g_addr_bits-1 downto 0);
		i_data		: in std_logic_vector(g_width-1 downto 0);
		o_data		: out std_logic_vector(g_width-1 downto 0));
end ram_l2_n7;

architecture rtl of ram_l2_n7 is
	type t_mem is array (0 to g_depth-1) of std_logic_vector(g_width-1 downto 0);
	signal r_mem : t_mem := ("1111111111000010", "0000000100011101", "1111010001001100", "1111111110010011", "0000000000000001", "0000000001100010", "0000110011101111", "0000001001010000", "0000000000011000", "0000000001001111", "1111111010101010", "1111111111100110", "1111111110110101", "0000101100101100", "0000101011001110", "0000000000111000", "0000110010110011", "0000000000001100", "0000000001011101", "1111111111101011", "1111011011111100", "1111111111111111", "0000000000101011", "1111100111111001", "0000001011010101", "1111111101011001", "0000000000010011", "1111001111011100", "0000000001100010", "0000000001100101" , others => (others => '0'));

begin
	p_ram : process(i_clk)
	begin
		if rising_edge(i_clk) then
			if (i_wr='1') then
				r_mem(to_integer(unsigned(i_addr))) <= i_data;
			end if;
			o_data <= r_mem(to_integer(unsigned(i_addr)));
		end if;	end process p_ram;end rtl;