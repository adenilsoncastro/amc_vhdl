library ieee;
 use ieee.std_logic_1164.all;
 use ieee.numeric_std.all;
 
 entity ram is
	generic(
		g_width 		: natural := 16;
		g_depth 		: natural := 863;
		g_addr_bits : natural := 10);
	
	port(
		i_clk			: in std_logic;
		i_wr			: in std_logic;
		i_addr		: in std_logic_vector(g_addr_bits-1 downto 0);
		i_data		: in std_logic_vector(g_width-1 downto 0);
		o_data		: out std_logic_vector(g_width-1 downto 0));
 end ram;
 
 architecture rtl of ram is
	type t_mem is array (0 to g_depth-1) of std_logic_vector(g_width-1 downto 0);
	signal r_mem : t_mem := 
	("0000000000000000","0000000000110001","1111111101100000","0000000000110100","1111111110101111",
	"0000000000101100","0000000001010100","0000000011110010","0000111111110110","1111111100100011",
	"0000001111011010","0000001011100100","1111100111000000","1111110110001101","0000000010111010",
	"0000110000101001","1111110100111011","0000101011111000","0000011010011010","0000111101111100",
	"0000001011110110","0000000100101110","0000111010111011","1111111110000011","1111001101101111",
	"1110001110011001","0000010100101000","0000010011010100","0000001101011101","0001010100010001",
	"0000000101010010","0000100101011001","1111110001010111","1111111110111011","0000001010110110",
	"0000000010100101","1111101110000011","1111111110101110","1101011000100111","0000011111110110",
	"1111001111110011","0000100100111100","1111110011001000","1111111101011100","1111101011011000",
	"0001001011101100","0001101101010101","0000001110110011","0001100010001100","0000001000110010",
	"0000000100100111","0000000111111110","1110110101010001","0001001010011011","1111111100011101",
	"1100111010000001","0000001000101011","1111111100110001","0000001000110110","1110111001101100",
	"0001001100111100","1111111001001001","1101000010110101","0000010010100100","1111111110000101",
	"1111101001001011","1111110000011000","1111110111110101","1111101010101101","1111100111001100",
	"1111110000000001","1111111000000011","0000010001011111","0000001011111001","0000000010001100",
	"0000011001010101","1111100001010000","1111110001101011","0000000100000101","0000001001001100",
	"0000110001001000","1110110011000100","0000010110011100","0010001011000100","0000001000110101",
	"0000000000101110","0000000110110001","1111000001011000","0001001111110100","1111111001111010",
	"1100111100111110","1111101010111011","0000000101110010","0000010111110010","1111110000001001",
	"0001000110111110","0000101111000011","0000111000011111","1111110101000001","1111111110101000",
	"1111100101010001","0001001001101001","0000110011111100","0000001011000010","0001110001100100",
	"1111101101111000","0000000101010000","0000011010010100","0000001001010010","0000001000011010",
	"0000010101101111","1101110100111101","0000001101000001","0000000100011000","0000011101101110",
	"1110110001000010","1110111001001010","1111101101001101","1110001000001011","0000000111000100",
	"0000000100001000","1111110000001110","0001010000011110","1111101011110000","1111011111100011",
	"0001101001110110","0000001110101001","0000000001011111","0000011101101100","1110111110100000",
	"1110011000000000","1111101011000010","1110011111111010","0000010101001010","0000000110110111",
	"1111011011101101","0000010000000010","1110101100111110","1111010111000000","1111000001110001",
	"0000010100011000","1111111111010010","1111100001001110","1111110001100011","1111110100110101",
	"1111101010101101","0000100000001011","0000010100000100","1111111010111001","1111100001110010",
	"1111110011010011","1111110110000111","1111101001110001","0000101100000000","0000001000010010",
	"1111111111010011","0000000000101000","1111000001111111","0001010000001100","1111110111100101",
	"1100110110101001","0000001011110111","0000000000010110","0000000010010000","1110111111011101",
	"0001010011101110","1111110000010010","1100111110100111","0000010100000011","0000000000101111",
	"1111100011100001","1111110001111110","1111110111100101","1111101010110000","0000110011001011",
	"1111111100000111","1111111011000000","0000001111101100","1110101010100110","0000100001001001",
	"0000011000011101","1110000011000100","0000010100111011","1111111110101111","1111100100000111",
	"1111110101001011","1111111001000011","1111101000100101","0001010110110100","1111101011111000",
	"1111111101100001","0000010111110010","0000001111000111","0000000101101100","0000010111000011",
	"1111001000000010","0000001000111100","0000001001101111","0000011110011100","1110110101101000",
	"1111001001000100","1111110101101111","1110010011001000","1111101011000011","1111111101110001",
	"0000001010011000","0000100011111011","0010000001101100","0000100100001100","0001001000011001",
	"0000000010000010","0000000011111010","1111101111011011","0001011111001000","1111100100010010",
	"1111100111010000","0001111111101100","0000010011111101","1111111111111101","1111100100011000",
	"1111110101110110","1111111000100100","1111101001010001","0001101011101001","0000010100101000",
	"1111111100110000","1111100010101110","1111110101001110","1111111001010011","1111101000011001",
	"0000011110011110","0000001101011001","1111111110000000","1111100000011011","0000111010011000",
	"1111100100000111","1111010101101100","1111111000011010","0000001011001010","1111111011000111",
	"0000011110110011","1110111000101000","1111000111111010","1111110001111100","1110010010010100",
	"1111110100010010","0000000000111001","1111100100001011","0001001010010011","0001000111001100",
	"0000001101001111","0001100110000010","1111110000111011","0000001000100111","0000100000100010",
	"0000100000101010","0000000111111101","1111110000111001","1111011111000111","0000100001000010",
	"1111101010100101","0000001101011100","1111111000110000","1111111000100010","0000000100000100",
	"1111111000100011","0000010100110011","0000000100001100","0000000100011101","0000100001100010",
	"0000100100011000","0000000110000000","0000000100001101","0000000011101001","1111111001100010",
	"1111111010001000","1111111011011101","1111111001111011","0000000101110111","0000000001111111",
	"0000001111000100","1111110101001101","0000000011011110","0000000001110010","1111110010100010",
	"0000000001010000","1111111101101011","1111111111111100","0000000010101001","1111111110000111",
	"1111111011011100","1111111011111010","1111110001010101","0000000010100101","0000001110100000",
	"0000000000000110","0000001101011000","0000001000011101","1111111100111100","1111111111010001",
	"0000000010100100","1111111111100001","1111111110000001","0000000010000110","1111111111110000",
	"1111111111011101","0000010011111000","1111110101011001","1111111011011010","1111111110000000",
	"1111111100111110","1111111011110010","0000010101001011","1111101100110101","0000001000001110",
	"0000011010100000","1111110100011011","1111101111011010","1111111101000010","1111111110001101",
	"0000010110111000","1111110000011000","0000010101001100","0001001010011110","1111111100100101",
	"1111000001001000","0000001000110110","1111100000011110","1111101111010101","1111111101001001",
	"0000000010010010","1111101111000011","1111101100001111","0000000010001100","1111110001110010",
	"0000000010000110","1111111110001100","1110111110101100","0000011100110111","0000001010110101",
	"1111111100100101","1111111111101000","1111110011110000","1110111111100101","0000110001011101",
	"1111111101101000","0000000000111010","1111111011100100","1111111011000111","1111010111000111",
	"0000000110011010","0000000000001001","1111111010000110","1111111110111111","1111111110011000",
	"0000010111111010","1111111111011111","0000000000100011","0000000000111010","1111111111101100",
	"1111001100000011","1111010011011110","1111111101010111","1111111110111010","1111010001101111",
	"0000000000010111","1111010100011100","0000101000000000","0000000000100100","1111111111000100",
	"1111111101011110","1111011001001110","1111001010111100","0000000010010010","1111111111110100",
	"0000000011101011","0000000011110111","0000000101111000","1111110011011000","1111110000010100",
	"1111101111010100","0000101001011010","0000000100100001","1111110100000010","0000000000110110",
	"0000001001010011","0000011000000011","1111111000111001","0000000111101011","1111111110010111",
	"0000000001111001","1111110100111101","1111110010000101","1111110101000000","1111111001010001",
	"1111110010001000","1111110011110101","1111110000010111","0000010010111000","1111110100110101",
	"0000000110100110","0000001111100011","1111101111100010","1111111001011111","0000000101111110",
	"1111110111100111","0000001011111110","0000000011011010","0000100011010101","0000010010111010",
	"0000010001101110","1111110011000110","0000001010100101","0000001111001001","0000010110101101",
	"0000111001101111","0000011100010101","0000001000100010","1111011010111101","1111101111000110",
	"1111011100011100","1111010000001010","1111110110101001","1111110111100001","0000010000101110",
	"0000000100101001","1111110101100101","0000010011101101","1111111001110000","0000000101111010",
	"1111100000100001","0001000111111001","1111101111000000","1111110101101001","1111110110010011",
	"1111100111000110","1111011110101010","0000101001011100","1111111011110111","0000000001101011",
	"0000011100011011","0000010110001101","0000000011111110","1111111011010001","1111111001000110",
	"0000011001101101","1111111110001010","1111111010110001","1111111110011100","0000000000110100",
	"1111110001100100","1111111101111111","0000000001110001","0000000000101101","0000000001111100",
	"0000010011111011","0000010001010110","0000000001010010","0000010001011010","0000000000110110",
	"1111111100100010","0000000110010001","0000000001010101","1111101000110111","0000000010101001",
	"0000000010011110","0000000100111001","0000000010010100","1111111100010000","0000000001011110",
	"1111111111100111","0000000011010101","0000000011011111","0000100101000011","1111111100011110",
	"1111111110011100","0000000001101110","1111111111010110","1111111111100101","1111101010000110",
	"0000000010000100","1111111110010000","1111111111110101","1111111111100100","0000101010000011",
	"0000101001100010","0000000001011001","0000000000001001","0000110000110011","0000000101100010",
	"0000101001101011","1111011000010001","0000000000011111","1111111111110001","1111111100101111",
	"0000100010001010","0000101001100110","0000000000010101","0000000000010011","0000000010101111",
	"1111111101001100","1111111111010110","1111111011000011","1111111100010001","1111011110110010",
	"0000000111101110","0000000001100011","1111111111101101","0000000000011010","0000000001100100",
	"0000011110000000","1111111110101111","1111111110110011","1111111111110101","1111111111000000",
	"1111001110111111","1111010000101101","1111111010111000","1111111110100110","1111001111100100",
	"1111111100110001","1111010000111011","0000101000100010","0000000010000001","0000000000001100",
	"0000000010111111","1111010110010100","1111010101110010","0000000001110011","0000000001110101",
	"1111111110010100","0000100000010011","1111000010100111","0000110011010001","0000110011100011",
	"1111101100010101","0000011001000101","1111111111110100","0000011111010001","0001000010011010",
	"1110010110010010","0000001011000010","0001011100010011","1110000111010101","0001000100111111",
	"1111000101111101","1111101100011001","1111110010010011","0000010010000000","0000010010100101",
	"1111101111000010","0001111001111010","1111110110011101","0000001111100010","0001111100011111",
	"0000001101001011","1101111010010011","1111110110010010","1111110001110101","1110010001000110",
	"0001101000010000","1110101110011111","1111110101001100","1111101101101001","1111100100101000",
	"1111100100000000","0000010110011100","1111101010111110","0000000011001100","1111110001110011",
	"1110000011111010","0000001011101000","1111111001100101","1111111001111011","0000101100101111",
	"0000010110100110","0001011110011000","0000001111010001","0000001101101011","1111101010110100",
	"1111110100100101","0000010001001011","1111001001010110","0000000100100101","1111110100111110",
	"1111111100100010","1111010010011110","0000101110011000","0000001010100101","0000001101101101",
	"0001111100010000","1111110101111000","1111111011001111","0000000100100110","1111111110000011",
	"0000000111100100","0000001010001110","0001000110100110","0000000111010111","1111111100001001",
	"0000001001111011","1111111101010011","1111111100001001","0000000111101000","0000000011101001",
	"0000000101110110","0000000001110101","0000000010110110","0000011101011011","0000010111111010",
	"0000000110011101","0000001000110101","0000001010111010","1111111111010011","0000010100100000",
	"1111110110011111","0000000101001001","1111111110100001","0000000100001011","0000001010011100",
	"0000100101110010","0000000011110010","0000000101001110","1111111011100110","1110100001101100",
	"0000000110111110","1111011001010010","1111100100001100","1111011011100101","1111101010111011",
	"1111001011010011","1111011011110010","0000100001001001","1111100100011001","1110011001010010",
	"0001011111001100","0001011100000100","1111111111101010","0000010110101010","0001010101001111",
	"1111001001110011","0000100010011000","1111111000111010","1111010100010110","0000011110001110",
	"1111010111011110","0000100011011001","0000011111110111","1111110101010101","1111011100101011",
	"1101110101010101","0010111100011011","1110100101010100","0000100011010111","1111101100000101",
	"1110101001010110","0000001111110011","0010000101011111","0000010000011111","1111101100100111",
	"1111101010010011","1111110101101100","0000011000100111","0000001001001011","1111101100101011",
	"1110001111010111","0000101101100000","1111110100001001","0000010110111101","0000100001011100",
	"1111100001111010","0000001110111100","1111110000101010","1111110000001111","0000001000111110",
	"0000001000010001","1111110011001100","0000000011111000","1111110100010011","0000000011001001",
	"0100010111010100","0000000001011001","0000000010000110","1111110110010110","1011001100111101",
	"0100011000010101","1111111101111001","1111111111101000","1100110010000100","0010010010101011",
	"1111111110001000","0000101101110111","1111100010000111","0000001101001101","0000110111111111",
	"0001001000100010","0010011111101011","1111110001100101","0000010100110011","0010100000100000",
	"1101111100100010","1111101111000101","0000011100011111","1111110010000011","0000010111011100",
	"1111110001100000","1111110100011101","0000100001100001","1111110111010111","1111101101000010",
	"0000001010100010","1111110101101100","0000000011100011","0000000000111000","0000011010100100",
	"0000010011010001","1111001011100111","1111001111011100","0000010100111001","0000100000101101",
	"0011100110000011","0000011011111100","1110101110000000","1111011001010101","0000100110111101",
	"0000000001010001","1111111001000110","1111000110100101","0001011101101100","1111100100100101",
	"1101101010110100","0000100111000101","0000011000010011","0000011001010110","0011000001000010",
	"0001011101010101","1111100010111110","0000011000000010","0000001010010001","1101010000110000",
	"1111100010000001","1111100010000001","0000001111110110","0001101011100001","1111011101000011",
	"1111111101010111","1111010001111011","1101101100110011","1111010001011100","1111111101111101",
	"1111111110101010","1111100011111111","0000101101110011","0000001000101101","1110001010010010",
	"1111101111010011","1111011011101101","1111110101111000","1111101000010101","0000111010001010",
	"0000001010110011","1111010001000100","0000010111010100","1111101001010011","1111011011101110",
	"0000110000011001","0000000111011001","1111110000000110","0001000001001110","0000000110101111",
	"1111111001110011","1110011011010110","1110011111001000","1111001110100000","0000001100110101",
	"0001101110001001","1110011000110101","1111011110110011","0000010110100010","0010000100100101",
	"1110111110100011","0001011000001111","0001111011010011","1110011111100110","1111111011101001",
	"1111110011111000","1111010010110001","0011000000011010","0000000101010111","1111111100010001",
	"0000001010111110","0000100000100100","0000000011010111","1110101101001011","0010000101101100",
	"0010101100111010","0000100001101001","1111111111001110","1111101110000110","1111010101000001",
	"1101001101011111","0010111010011010","1110110100000001","1111000111111010","0011010110100101",
	"0010011111110001","1111111100111100","1110110001101101","0000011110001101","0000110011001010",
	"0000011101110011","1110111000101110","0000101101110010","1110010010010010","1111100011101011",
	"1110100010111101","1110010101011001","0010001001111111","0000011000100111","0000011111011011",
	"1110101011010000","1111000010011100","0001001000111101","0001010000111000","0011101111110010",
	"1111111101010101","0000101010000100","0000110111110111","1111110111100100","1110001101101100",
	"0000111011101010","0000010001011110","0001001110101001","0000011010010110","0001101010101101",
	"1111111101010000","0000101110101101","1111100001000001","0000110101011001","1101000000100010",
	"0000110101010011","0000010010000001","1111010110111000","1111000100101010","1110001100010001",
	"0000110111011010","1111101001111101","0000010101111000","0010111111110100","1110010100011011",
	"1111101110110100","0000101010110000","0000000100001101","1110000100001010","0111111111111111",
	"1110010000101011","1111101001110101","0000000111000101","1111001110101011","0001110001000111",
	"0000001000111000","1101010011010101","0010101000100100");
	
 begin
	p_ram : process(i_clk)
	begin
		if rising_edge(i_clk) then
			if (i_wr='1') then
				r_mem(to_integer(unsigned(i_addr))) <= i_data;
			end if;
			o_data <= r_mem(to_integer(unsigned(i_addr)));
		end if;
	end process p_ram; 
 end rtl;