-- megafunction wizard: %ALTMULT_ACCUM (MAC)%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altmult_accum 

-- ============================================================
-- File Name: mac_alt.vhd
-- Megafunction Name(s):
-- 			altmult_accum
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2020  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY mac_alt IS
	PORT
	(
		clock0		: IN STD_LOGIC  := '1';
		dataa		: IN STD_LOGIC_VECTOR (7 DOWNTO 0) :=  (OTHERS => '0');
		datab		: IN STD_LOGIC_VECTOR (7 DOWNTO 0) :=  (OTHERS => '0');
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END mac_alt;


ARCHITECTURE SYN OF mac_alt IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);



	COMPONENT altmult_accum
	GENERIC (
		accum_direction		: STRING;
		addnsub_aclr		: STRING;
		addnsub_pipeline_aclr		: STRING;
		addnsub_pipeline_reg		: STRING;
		addnsub_reg		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a		: STRING;
		input_aclr_b		: STRING;
		input_reg_a		: STRING;
		input_reg_b		: STRING;
		input_source_a		: STRING;
		input_source_b		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier_aclr		: STRING;
		multiplier_reg		: STRING;
		output_aclr		: STRING;
		output_reg		: STRING;
		port_addnsub		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		sign_aclr_a		: STRING;
		sign_aclr_b		: STRING;
		sign_pipeline_aclr_a		: STRING;
		sign_pipeline_aclr_b		: STRING;
		sign_pipeline_reg_a		: STRING;
		sign_pipeline_reg_b		: STRING;
		sign_reg_a		: STRING;
		sign_reg_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			clock0	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(15 DOWNTO 0);

	altmult_accum_component : altmult_accum
	GENERIC MAP (
		accum_direction => "ADD",
		addnsub_aclr => "UNUSED",
		addnsub_pipeline_aclr => "UNUSED",
		addnsub_pipeline_reg => "CLOCK0",
		addnsub_reg => "CLOCK0",
		dedicated_multiplier_circuitry => "YES",
		input_aclr_a => "UNUSED",
		input_aclr_b => "UNUSED",
		input_reg_a => "CLOCK0",
		input_reg_b => "CLOCK0",
		input_source_a => "DATAA",
		input_source_b => "DATAB",
		intended_device_family => "Cyclone IV E",
		lpm_type => "altmult_accum",
		multiplier_aclr => "UNUSED",
		multiplier_reg => "CLOCK0",
		output_aclr => "UNUSED",
		output_reg => "CLOCK0",
		port_addnsub => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "SIGNED",
		representation_b => "SIGNED",
		sign_aclr_a => "UNUSED",
		sign_aclr_b => "UNUSED",
		sign_pipeline_aclr_a => "UNUSED",
		sign_pipeline_aclr_b => "UNUSED",
		sign_pipeline_reg_a => "CLOCK0",
		sign_pipeline_reg_b => "CLOCK0",
		sign_reg_a => "CLOCK0",
		sign_reg_b => "CLOCK0",
		width_a => 8,
		width_b => 8,
		width_result => 16
	)
	PORT MAP (
		clock0 => clock0,
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ACCUM_SLOAD NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR NUMERIC "3"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_ACLR NUMERIC "3"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG NUMERIC "1"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG_INDEX NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_REG NUMERIC "1"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_REG_INDEX NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_ACLR NUMERIC "3"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_ACLR NUMERIC "3"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_REG NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_REG NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
-- Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "0"
-- Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "0"
-- Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: EXTRA_MULTIPLIER_LATENCY NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_MAC STRING "1"
-- Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "1"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: MULT_LATENCY NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "1"
-- Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "1"
-- Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "1"
-- Retrieval info: PRIVATE: NUM_MULT STRING "1"
-- Retrieval info: PRIVATE: OP1 STRING "Add"
-- Retrieval info: PRIVATE: OP3 STRING "Add"
-- Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
-- Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: OVERFLOW NUMERIC "0"
-- Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: REG_OUT NUMERIC "1"
-- Retrieval info: PRIVATE: RNFORMAT STRING "16"
-- Retrieval info: PRIVATE: RQFORMAT STRING "Q1.30"
-- Retrieval info: PRIVATE: RTS_WIDTH STRING "16"
-- Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
-- Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
-- Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
-- Retrieval info: PRIVATE: SCANOUTA NUMERIC "0"
-- Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
-- Retrieval info: PRIVATE: SIGNA STRING "SIGNED"
-- Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNA_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNB STRING "SIGNED"
-- Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNB_REG STRING "1"
-- Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIDTHA STRING "8"
-- Retrieval info: PRIVATE: WIDTHB STRING "8"
-- Retrieval info: PRIVATE: WIDTH_UPPER_DATA NUMERIC "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ACCUM_DIRECTION STRING "ADD"
-- Retrieval info: CONSTANT: ADDNSUB_ACLR STRING "UNUSED"
-- Retrieval info: CONSTANT: ADDNSUB_PIPELINE_ACLR STRING "UNUSED"
-- Retrieval info: CONSTANT: ADDNSUB_PIPELINE_REG STRING "CLOCK0"
-- Retrieval info: CONSTANT: ADDNSUB_REG STRING "CLOCK0"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "YES"
-- Retrieval info: CONSTANT: INPUT_ACLR_A STRING "UNUSED"
-- Retrieval info: CONSTANT: INPUT_ACLR_B STRING "UNUSED"
-- Retrieval info: CONSTANT: INPUT_REG_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A STRING "DATAA"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B STRING "DATAB"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_accum"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR STRING "UNUSED"
-- Retrieval info: CONSTANT: MULTIPLIER_REG STRING "CLOCK0"
-- Retrieval info: CONSTANT: OUTPUT_ACLR STRING "UNUSED"
-- Retrieval info: CONSTANT: OUTPUT_REG STRING "CLOCK0"
-- Retrieval info: CONSTANT: PORT_ADDNSUB STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
-- Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
-- Retrieval info: CONSTANT: SIGN_ACLR_A STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGN_ACLR_B STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGN_PIPELINE_ACLR_A STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGN_PIPELINE_ACLR_B STRING "UNUSED"
-- Retrieval info: CONSTANT: SIGN_PIPELINE_REG_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGN_PIPELINE_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGN_REG_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGN_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "16"
-- Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
-- Retrieval info: USED_PORT: dataa 0 0 8 0 INPUT GND "dataa[7..0]"
-- Retrieval info: USED_PORT: datab 0 0 8 0 INPUT GND "datab[7..0]"
-- Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT GND "result[15..0]"
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 8 0 dataa 0 0 8 0
-- Retrieval info: CONNECT: @datab 0 0 8 0 datab 0 0 8 0
-- Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
-- Retrieval info: LIB_FILE: altera_mf
